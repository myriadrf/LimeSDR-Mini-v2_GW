// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.12.1.454
// Netlist written on Sun Jan 23 21:09:16 2022
//
// Verilog Description of module top
//

module top (REF_CLK, USER_BUTTON, LED_R, LED_G, LED_B, IO_SCK, IO_MOSI, 
            IO_MISO, IO_0);   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(21[8:11])
    input REF_CLK;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    input USER_BUTTON;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(24[7:18])
    output LED_R;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(25[7:12])
    output LED_G;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(26[3:8])
    output LED_B;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(27[3:8])
    output IO_SCK;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(28[3:9])
    output IO_MOSI;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(29[3:10])
    output IO_MISO;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(30[3:10])
    output IO_0;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(31[3:7])
    
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(59[8:24])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(59[8:24])
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire IO_SCK_c /* synthesis is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(28[3:9])
    wire sclk_N_5010 /* synthesis is_inv_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(57[11:19])
    
    wire USER_BUTTON_c, LED_R_c_0, LED_G_c_0, LED_B_c_0, IO_MOSI_c, 
        IO_MISO_c, IO_0_c_0, inst1_FIFOif_rd, inst1_FIFOof_wr, inst1_FIFOfifo_rst;
    wire [15:0]\from_fpgacfg.phase_reg_sel ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    wire [4:0]\from_fpgacfg.clk_ind ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    wire [4:0]\from_fpgacfg.cnt_ind ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    
    wire \inst2_from_fpgacfg.load_phase_reg ;
    wire [15:0]\from_fpgacfg.drct_clk_en ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    wire [15:0]\from_fpgacfg.ch_en ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    wire [1:0]\from_fpgacfg.smpl_width ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    
    wire \inst2_from_fpgacfg.mode , \inst2_from_fpgacfg.ddr_en , \inst2_from_fpgacfg.trxiq_pulse , 
        \inst2_from_fpgacfg.mimo_int_en , \inst2_from_fpgacfg.synch_dis , 
        \inst2_from_fpgacfg.synch_mode , \inst2_from_fpgacfg.smpl_nr_clr , 
        \inst2_from_fpgacfg.txpct_loss_clr , \inst2_from_fpgacfg.rx_en , 
        \inst2_from_fpgacfg.tx_en , \inst2_from_fpgacfg.rx_ptrn_en , \inst2_from_fpgacfg.tx_ptrn_en , 
        \inst2_from_fpgacfg.tx_cnt_en ;
    wire [15:0]\from_fpgacfg.wfm_ch_en ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    wire [15:0]n33_adj_6951;
    
    wire \inst2_from_fpgacfg.wfm_load ;
    wire [1:0]\from_fpgacfg.wfm_smpl_width ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    wire [15:0]\from_fpgacfg.SPI_SS ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    
    wire \inst2_from_fpgacfg.LMS1_SS , \inst2_from_fpgacfg.LMS1_RESET , 
        \inst2_from_fpgacfg.LMS1_CORE_LDO_EN , \inst2_from_fpgacfg.LMS1_TXNRX1 , 
        \inst2_from_fpgacfg.LMS1_TXNRX2 , \inst2_from_fpgacfg.LMS1_TXEN , 
        \inst2_from_fpgacfg.LMS1_RXEN ;
    wire [15:0]\from_fpgacfg.GPIO ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    wire [2:0]\from_fpgacfg.FPGA_LED1_CTRL ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    wire [2:0]\from_fpgacfg.FPGA_LED2_CTRL ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    wire [2:0]\from_fpgacfg.FX3_LED_CTRL ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    wire [3:0]\from_fpgacfg.CLK_ENA ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    wire [31:0]\from_fpgacfg.sync_pulse_period ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    wire [15:0]\from_fpgacfg.sync_size ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    wire [15:0]\from_fpgacfg.txant_pre ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    wire [15:0]\from_fpgacfg.txant_post ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(40[7:19])
    wire [31:0]inst3_Q;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(62[8:15])
    
    wire inst3_Empty, inst3_Full, n3;
    wire [15:0]inst_reg;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(51[11:19])
    
    wire n2, n41299, n41298;
    wire [31:0]SHAREDBUS_ADR_I;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(361[13:28])
    wire [31:0]SHAREDBUS_DAT_I;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(362[13:28])
    wire [31:0]LM32I_ADR_O;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(376[13:24])
    
    wire locked_N_493;
    wire [31:0]LM32D_ADR_O;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(389[13:24])
    
    wire n45106, n45105;
    wire [1:0]selected;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(244[15:23])
    wire [2:0]LM32D_CTI_O;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(397[12:23])
    
    wire LM32D_CYC_O, n145, n41292;
    wire [2:0]counter;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(465[11:18])
    
    wire n37509, n37508, n37507, n37506, REF_CLK_c_enable_1424, n6518, 
        n37505, n37504, n37503, n37502, n37501, n37500, n37499, 
        n37498, n37497, n37496, n37495, n5386, n10865, n2023, 
        n6439, n6781, n6589, n148, n85, n6512, n142, n139, n151, 
        n45076, n45103, n45101, n45099, n6604, n109, n133, n6502, 
        n136, n82, n130, n19822, n103, n79, n6584;
    wire [14:0]\genblk1.pmi_address ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(242[31:42])
    
    wire n6640;
    wire [12:0]\genblk1.read_address ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(243[31:43])
    wire [12:0]\genblk1.write_address ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(243[45:58])
    wire [2:0]\genblk1.state ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(255[13:18])
    
    wire n27508, n3486, n3485, n3432, n6609, n5085;
    wire [0:0]PIO_DATAI_adj_6643;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/gpio/rtl/verilog/gpio.v(146[27:36])
    
    wire n27507, n36339, n124, n6429, n27506, rx_shift_data_31__N_4339, 
        n6624, n34242, n27505, n41263, n37;
    wire [31:2]branch_target_d;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(397[21:36])
    
    wire n36;
    wire [4:0]write_idx_w;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(476[25:36])
    wire [31:0]w_result;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(521[22:30])
    wire [31:0]operand_1_x;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(524[22:33])
    wire [31:0]operand_m;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(526[22:31])
    wire [31:0]adder_result_x;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(559[23:37])
    
    wire n34;
    wire [31:0]shifter_result_m;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(583[23:39])
    wire [31:2]pc_f;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(631[21:25])
    wire [31:2]pc_d;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(632[21:25])
    
    wire dcache_refill_request, dc_re, n27503, n6599, n6515, n27502, 
        n32312, n76, n73, n64, n70, n67, n6764, n6763, n6762, 
        n6761, n6760, n100, n6424, n6619, n27501, REF_CLK_c_enable_164, 
        n94, n88, n91, n118, n121, n97, n27500, n27499, n27498, 
        n27497, n127, n27496, n27495, n27494, n30231, n27493, 
        dcache_select_x;
    wire [31:0]dcache_refill_address;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(254[23:44])
    wire [2:0]next_cycle_type_adj_6725;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(257[24:39])
    
    wire n6759, n6614, n27492, n27491, n27490;
    wire [31:0]d_adr_o_31__N_2278;
    
    wire n27489, n106, n34_adj_6597, n37_adj_6598, n6758, n27488, 
        n27487, direction_m;
    wire [31:0]left_shift_result;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(93[22:39])
    
    wire n40, n43, n46, n49, n52, n55, n58, n61, n64_adj_6599, 
        n67_adj_6600, n112, n70_adj_6601, n73_adj_6602, n27486, n76_adj_6603;
    wire [31:0]p;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(132[22:23])
    wire [31:0]a;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(133[22:23])
    wire [31:0]b;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(134[22:23])
    wire [32:0]t;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(136[13:14])
    
    wire n6757, n6756, n27485, n27483, n115, bie, n35448, n27482, 
        n27481, n7676, n7675, n7674, n7673, n7672, n7671, n7670, 
        n7669, n7668, n7667, n7666, n7665, n7664, n7663, n7662, 
        n7661, n7660, n35647, n27480, n7659, n7658, n7657, n7656, 
        n27479, n7655, n7654, n6434, n27478, n27477, n8, n27476, 
        n27475, n6038, bie_N_3274, n29830, n6034, n7653, n7652, 
        n7651, n7650, n7649, n7648, n7647, n7646, n7645, n7644, 
        n7643, n7642, n7641, n7640, n7639, n7638, n7637, n7636, 
        n7635, n7634, n7633, n7632, n7631, n7630, n7629, n7628, 
        n7627, n7626, n7625, n7624, n7623, n7622, n10452, n6637, 
        n27474, n27473, n27472, n7621, n7620, n7619, n7618, n7617, 
        n7616, n7615, n7614, n7613, n7611, n7610, n7608, n7607, 
        n7606, n7605, n7604, n7603;
    wire [8:0]flush_set;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(200[30:39])
    
    wire n7602, n7601, n27471, n27470;
    wire [8:0]flush_set_8__N_1953;
    
    wire n6755, n6754, n6753, n6629, n7600, n7599, n7598, n7597, 
        n7596, n7595, n7594, n7593, n7592, n7591, n7590, n7589, 
        n7588, n7587, n7586, n7585, n7584, n7583, n7582, n7581, 
        n7580, n7579, n7578, n7577, n7576, n7575, n7574, n7573, 
        n7572, n7571, n6642, n7570, n7569, n7568, n7567, n7566;
    wire [8:0]tmem_write_address_adj_6794;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(180[31:49])
    wire [10:0]dmem_write_address_adj_6796;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(182[31:49])
    wire [2:0]state_adj_6798;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(186[26:31])
    wire [8:0]flush_set_adj_6801;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(195[30:39])
    wire [8:0]flush_set_8__N_2513;
    
    wire n6752, n6751, n6750, n7565, n7564, n7563, n7562, n7561, 
        n7560, n7559, n7558, n7557, n7556, n7555, n7554, n7553, 
        n7552, n7551, n7550, n7549, n7548, n7547, n7546, n7545, 
        n6645, n6648, n6749, n36319, n27469, n12428, n27468, n27467, 
        n27466, n6574, n6594, n36321, n36330, n6579, n36329, n3700, 
        n27465, n27464, n27463, n36325, n36336, n36337, n11843, 
        n31279, n27462, n36326, n27460, n36320, n36340, n10587, 
        n10589, n10591, n10593, n10595, n41191, n27459, n27458, 
        n36322, n27457, n27456, n27455, n36332, n36331, n36328, 
        n27454, n36335, n36338, n29, REF_CLK_c_enable_176, REF_CLK_c_enable_161, 
        n10585, n27453, n27452, n27451, n27450, n27449, n27448, 
        n27447, n35006, n17816, n34966, n27446, n27445, n27444, 
        n45086, n38965, n38964, n27443, n27442, n38963, n41434, 
        n41432, n41430, n34926, n27441, n36323, n27440, n41425, 
        n27439, REF_CLK_c_enable_1606, n27438, n36324, n36333, REF_CLK_c_enable_132, 
        n41405, REF_CLK_c_enable_158, n41401, REF_CLK_c_enable_177, 
        n41394, n41390, n36334, n41496, n41380, n41379, n41495, 
        n27437, n20000, n41359, n41358, n37240, n37239, n37238, 
        n37237, n37236, n37235, n37234, n37233, n37232, n37231, 
        n37230, n37229, n37228, n37227, n41357, n41356, n41355, 
        n37190, n37189, n37188, n37187, n37186, n37185, n37184, 
        n37183, n37182, n37181, n37180, n37179, n37178, n37177, 
        n37176, n41354, n41353, n41352, n41351, n41350, n41347, 
        n41346, n41344, n41343, n41342, n41341, n41340, n41339, 
        n41338, n41337, n41336, n41335, n41334, n41333, n41332, 
        n41331, n41330, n41329, n41328, n41325, n41321, n41310, 
        n41303, REF_CLK_c_enable_1453, n45179, n41301, n41300;
    
    VHI i2 (.Z(VCC_net));
    LUT4 i2744_4_lut (.A(n6512), .B(n37190), .C(n6515), .D(n41352), 
         .Z(n6518)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i2744_4_lut.init = 16'hc088;
    fpgacfg inst2 (.sclk_N_5010(sclk_N_5010), .n41434(n41434), .VCC_net(VCC_net), 
            .\from_fpgacfg.wfm_ch_en ({\from_fpgacfg.wfm_ch_en }), .REF_CLK_c(REF_CLK_c), 
            .\from_fpgacfg.CLK_ENA ({\from_fpgacfg.CLK_ENA }), .IO_MOSI_c(IO_MOSI_c), 
            .\from_fpgacfg.FX3_LED_CTRL ({\from_fpgacfg.FX3_LED_CTRL }), .\from_fpgacfg.FPGA_LED1_CTRL ({\from_fpgacfg.FPGA_LED1_CTRL }), 
            .\from_fpgacfg.GPIO ({\from_fpgacfg.GPIO }), .\from_fpgacfg.txant_post ({\from_fpgacfg.txant_post }), 
            .\from_fpgacfg.txant_pre ({\from_fpgacfg.txant_pre }), .\from_fpgacfg.sync_size ({\from_fpgacfg.sync_size }), 
            .\inst2_from_fpgacfg.wfm_smpl_width[0] (\from_fpgacfg.wfm_smpl_width [0]), 
            .\inst2_from_fpgacfg.rx_en (\inst2_from_fpgacfg.rx_en ), .\inst2_from_fpgacfg.smpl_nr_clr (\inst2_from_fpgacfg.smpl_nr_clr ), 
            .\from_fpgacfg.smpl_width ({\from_fpgacfg.smpl_width }), .\from_fpgacfg.ch_en ({\from_fpgacfg.ch_en }), 
            .\from_fpgacfg.clk_ind ({\from_fpgacfg.clk_ind }), .\from_fpgacfg.drct_clk_en ({\from_fpgacfg.drct_clk_en }), 
            .\from_fpgacfg.phase_reg_sel ({\from_fpgacfg.phase_reg_sel }), 
            .IO_0_c_0(IO_0_c_0), .\from_fpgacfg.SPI_SS ({\from_fpgacfg.SPI_SS }), 
            .\inst2_from_fpgacfg.load_phase_reg (\inst2_from_fpgacfg.load_phase_reg ), 
            .\inst2_from_fpgacfg.synch_mode (\inst2_from_fpgacfg.synch_mode ), 
            .\inst2_from_fpgacfg.tx_cnt_en (\inst2_from_fpgacfg.tx_cnt_en ), 
            .\from_fpgacfg.sync_pulse_period ({\from_fpgacfg.sync_pulse_period }), 
            .\inst2_from_fpgacfg.wfm_load (\inst2_from_fpgacfg.wfm_load ), 
            .\inst2_from_fpgacfg.wfm_play (n33_adj_6951[1]), .REF_CLK_c_enable_1424(REF_CLK_c_enable_1424), 
            .\inst2_from_fpgacfg.LMS1_RXEN (\inst2_from_fpgacfg.LMS1_RXEN ), 
            .\inst2_from_fpgacfg.LMS1_TXEN (\inst2_from_fpgacfg.LMS1_TXEN ), 
            .\inst2_from_fpgacfg.LMS1_TXNRX2 (\inst2_from_fpgacfg.LMS1_TXNRX2 ), 
            .\inst2_from_fpgacfg.LMS1_TXNRX1 (\inst2_from_fpgacfg.LMS1_TXNRX1 ), 
            .\inst2_from_fpgacfg.LMS1_CORE_LDO_EN (\inst2_from_fpgacfg.LMS1_CORE_LDO_EN ), 
            .\inst2_from_fpgacfg.LMS1_RESET (\inst2_from_fpgacfg.LMS1_RESET ), 
            .\from_fpgacfg.FPGA_LED2_CTRL ({\from_fpgacfg.FPGA_LED2_CTRL }), 
            .\inst2_from_fpgacfg.LMS1_SS (\inst2_from_fpgacfg.LMS1_SS ), .\inst2_from_fpgacfg.tx_en (\inst2_from_fpgacfg.tx_en ), 
            .\inst2_from_fpgacfg.rx_ptrn_en (\inst2_from_fpgacfg.rx_ptrn_en ), 
            .\inst2_from_fpgacfg.tx_ptrn_en (\inst2_from_fpgacfg.tx_ptrn_en ), 
            .\inst2_from_fpgacfg.txpct_loss_clr (\inst2_from_fpgacfg.txpct_loss_clr ), 
            .\inst2_from_fpgacfg.mode (\inst2_from_fpgacfg.mode ), .\inst2_from_fpgacfg.ddr_en (\inst2_from_fpgacfg.ddr_en ), 
            .\inst2_from_fpgacfg.trxiq_pulse (\inst2_from_fpgacfg.trxiq_pulse ), 
            .\inst2_from_fpgacfg.mimo_int_en (\inst2_from_fpgacfg.mimo_int_en ), 
            .\inst2_from_fpgacfg.synch_dis (\inst2_from_fpgacfg.synch_dis ), 
            .\from_fpgacfg.cnt_ind ({\from_fpgacfg.cnt_ind }), .n41191(n41191), 
            .\inst_reg[15] (inst_reg[15]), .REF_CLK_c_enable_1453(REF_CLK_c_enable_1453), 
            .n45086(n45086), .n10865(n10865), .n2023(n2023), .rx_shift_data_31__N_4339(rx_shift_data_31__N_4339), 
            .IO_MISO_c(IO_MISO_c), .n45179(n45179), .n35448(n35448), .USER_BUTTON_c(USER_BUTTON_c));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(110[9:28])
    CCU2C _add_1_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(b[0]), .B1(a[31]), .C1(GND_net), .D1(VCC_net), .COUT(n27445), 
          .S1(t[0]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam _add_1_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_add_4_2.INJECT1_1 = "NO";
    FD1P3DX creset_2683 (.D(n36319), .SP(REF_CLK_c_enable_161), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n6439));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_2683.GSR = "ENABLED";
    CCU2C add_22479_17 (.A0(adder_result_x[31]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27444), .S1(dcache_select_x));
    defparam add_22479_17.INIT0 = 16'h5555;
    defparam add_22479_17.INIT1 = 16'h0000;
    defparam add_22479_17.INJECT1_0 = "NO";
    defparam add_22479_17.INJECT1_1 = "NO";
    FD1P3DX creset_2675 (.D(n36320), .SP(REF_CLK_c_enable_176), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n6429));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_2675.GSR = "ENABLED";
    DPR16X4C n65110 (.DI0(n41425), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
            .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n6637), .RAD0(n41350), 
            .RAD1(n41354), .RAD2(n41351), .RAD3(n41353), .DO0(n6512));
    defparam n65110.initval = "0x0000000000000000";
    DPR16X4C n66440 (.DI0(write_idx_w[4]), .DI1(GND_net), .DI2(GND_net), 
            .DI3(GND_net), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n6640), .RAD0(n41355), .RAD1(n41358), .RAD2(n41359), 
            .RAD3(n41356), .DO0(n6645));
    defparam n66440.initval = "0x0000000000000000";
    FD1P3DX creset_2671 (.D(n36321), .SP(REF_CLK_c_enable_176), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n6424));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_2671.GSR = "ENABLED";
    CCU2C add_22479_7 (.A0(adder_result_x[21]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(adder_result_x[22]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n27439), .COUT(n27440));
    defparam add_22479_7.INIT0 = 16'h5555;
    defparam add_22479_7.INIT1 = 16'h5555;
    defparam add_22479_7.INJECT1_0 = "NO";
    defparam add_22479_7.INJECT1_1 = "NO";
    DPR16X4C registers0 (.DI0(w_result[28]), .DI1(w_result[29]), .DI2(w_result[30]), 
            .DI3(w_result[31]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n7611), .RAD0(n41350), .RAD1(n41354), .RAD2(n41351), 
            .RAD3(n41353), .DO0(n7605), .DO1(n7606), .DO2(n7607), .DO3(n7608));
    defparam registers0.initval = "0x0000000000000000";
    CCU2C add_22479_9 (.A0(adder_result_x[23]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(adder_result_x[24]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n27440), .COUT(n27441));
    defparam add_22479_9.INIT0 = 16'h5555;
    defparam add_22479_9.INIT1 = 16'h5555;
    defparam add_22479_9.INJECT1_0 = "NO";
    defparam add_22479_9.INJECT1_1 = "NO";
    DPR16X4C registers_d01 (.DI0(w_result[28]), .DI1(w_result[29]), .DI2(w_result[30]), 
            .DI3(w_result[31]), .WAD0(n45103), .WAD1(n45099), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n7610), .RAD0(n41355), 
            .RAD1(n41358), .RAD2(n41359), .RAD3(n41356), .DO0(n7641), 
            .DO1(n7642), .DO2(n7643), .DO3(n7644));
    defparam registers_d01.initval = "0x0000000000000000";
    DPR16X4C registers15 (.DI0(w_result[0]), .DI1(w_result[1]), .DI2(w_result[2]), 
            .DI3(w_result[3]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n7611), .RAD0(n41350), .RAD1(n41354), .RAD2(n41351), 
            .RAD3(n41353), .DO0(n7577), .DO1(n7578), .DO2(n7579), .DO3(n7580));
    defparam registers15.initval = "0x0000000000000000";
    DPR16X4C registers_d00 (.DI0(w_result[28]), .DI1(w_result[29]), .DI2(w_result[30]), 
            .DI3(w_result[31]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n7611), .RAD0(n41355), .RAD1(n41358), .RAD2(n41359), 
            .RAD3(n41356), .DO0(n7673), .DO1(n7674), .DO2(n7675), .DO3(n7676));
    defparam registers_d00.initval = "0x0000000000000000";
    DPR16X4C registers14 (.DI0(w_result[4]), .DI1(w_result[5]), .DI2(w_result[6]), 
            .DI3(w_result[7]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n7611), .RAD0(n41350), .RAD1(n41354), .RAD2(n41351), 
            .RAD3(n41353), .DO0(n7581), .DO1(n7582), .DO2(n7583), .DO3(n7584));
    defparam registers14.initval = "0x0000000000000000";
    DPR16X4C registers13 (.DI0(w_result[8]), .DI1(w_result[9]), .DI2(w_result[10]), 
            .DI3(w_result[11]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n7611), .RAD0(n41350), .RAD1(n41354), .RAD2(n41351), 
            .RAD3(n41353), .DO0(n7585), .DO1(n7586), .DO2(n7587), .DO3(n7588));
    defparam registers13.initval = "0x0000000000000000";
    DPR16X4C registers12 (.DI0(w_result[12]), .DI1(w_result[13]), .DI2(w_result[14]), 
            .DI3(w_result[15]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n7611), .RAD0(n41350), .RAD1(n41354), .RAD2(n41351), 
            .RAD3(n41353), .DO0(n7589), .DO1(n7590), .DO2(n7591), .DO3(n7592));
    defparam registers12.initval = "0x0000000000000000";
    DPR16X4C registers11 (.DI0(w_result[16]), .DI1(w_result[17]), .DI2(w_result[18]), 
            .DI3(w_result[19]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n7611), .RAD0(n41350), .RAD1(n41354), .RAD2(n41351), 
            .RAD3(n41353), .DO0(n7593), .DO1(n7594), .DO2(n7595), .DO3(n7596));
    defparam registers11.initval = "0x0000000000000000";
    DPR16X4C registers10 (.DI0(w_result[20]), .DI1(w_result[21]), .DI2(w_result[22]), 
            .DI3(w_result[23]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n7611), .RAD0(n41350), .RAD1(n41354), .RAD2(n41351), 
            .RAD3(n41353), .DO0(n7597), .DO1(n7598), .DO2(n7599), .DO3(n7600));
    defparam registers10.initval = "0x0000000000000000";
    DPR16X4C registers9 (.DI0(w_result[24]), .DI1(w_result[25]), .DI2(w_result[26]), 
            .DI3(w_result[27]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n7611), .RAD0(n41350), .RAD1(n41354), .RAD2(n41351), 
            .RAD3(n41353), .DO0(n7601), .DO1(n7602), .DO2(n7603), .DO3(n7604));
    defparam registers9.initval = "0x0000000000000000";
    DPR16X4C registers8 (.DI0(w_result[0]), .DI1(w_result[1]), .DI2(w_result[2]), 
            .DI3(w_result[3]), .WAD0(n45103), .WAD1(n45099), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n7610), .RAD0(n41350), 
            .RAD1(n41354), .RAD2(n41351), .RAD3(n41353), .DO0(n7545), 
            .DO1(n7546), .DO2(n7547), .DO3(n7548));
    defparam registers8.initval = "0x0000000000000000";
    DPR16X4C registers7 (.DI0(w_result[4]), .DI1(w_result[5]), .DI2(w_result[6]), 
            .DI3(w_result[7]), .WAD0(n45103), .WAD1(n45099), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n7610), .RAD0(n41350), 
            .RAD1(n41354), .RAD2(n41351), .RAD3(n41353), .DO0(n7549), 
            .DO1(n7550), .DO2(n7551), .DO3(n7552));
    defparam registers7.initval = "0x0000000000000000";
    DPR16X4C registers6 (.DI0(w_result[8]), .DI1(w_result[9]), .DI2(w_result[10]), 
            .DI3(w_result[11]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n7610), .RAD0(n41350), .RAD1(n41354), .RAD2(n41351), 
            .RAD3(n41353), .DO0(n7553), .DO1(n7554), .DO2(n7555), .DO3(n7556));
    defparam registers6.initval = "0x0000000000000000";
    DPR16X4C registers5 (.DI0(w_result[12]), .DI1(w_result[13]), .DI2(w_result[14]), 
            .DI3(w_result[15]), .WAD0(n45103), .WAD1(n45099), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n7610), .RAD0(n41350), 
            .RAD1(n41354), .RAD2(n41351), .RAD3(n41353), .DO0(n7557), 
            .DO1(n7558), .DO2(n7559), .DO3(n7560));
    defparam registers5.initval = "0x0000000000000000";
    DPR16X4C registers4 (.DI0(w_result[16]), .DI1(w_result[17]), .DI2(w_result[18]), 
            .DI3(w_result[19]), .WAD0(n45103), .WAD1(n45099), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n7610), .RAD0(n41350), 
            .RAD1(n41354), .RAD2(n41351), .RAD3(n41353), .DO0(n7561), 
            .DO1(n7562), .DO2(n7563), .DO3(n7564));
    defparam registers4.initval = "0x0000000000000000";
    DPR16X4C registers3 (.DI0(w_result[20]), .DI1(w_result[21]), .DI2(w_result[22]), 
            .DI3(w_result[23]), .WAD0(n45103), .WAD1(n45099), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n7610), .RAD0(n41350), 
            .RAD1(n41354), .RAD2(n41351), .RAD3(n41353), .DO0(n7565), 
            .DO1(n7566), .DO2(n7567), .DO3(n7568));
    defparam registers3.initval = "0x0000000000000000";
    CCU2C add_22479_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(adder_result_x[16]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n27437));
    defparam add_22479_1.INIT0 = 16'h0000;
    defparam add_22479_1.INIT1 = 16'haaaf;
    defparam add_22479_1.INJECT1_0 = "NO";
    defparam add_22479_1.INJECT1_1 = "NO";
    FD1P3DX creset (.D(n36322), .SP(REF_CLK_c_enable_161), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n6629));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset.GSR = "ENABLED";
    FD1P3DX creset_2807 (.D(n36323), .SP(REF_CLK_c_enable_132), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n6624));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_2807.GSR = "ENABLED";
    FD1P3DX creset_2803 (.D(n36324), .SP(REF_CLK_c_enable_132), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n6619));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_2803.GSR = "ENABLED";
    GSR GSR_INST (.GSR(VCC_net));
    FD1P3DX creset_2799 (.D(n36325), .SP(REF_CLK_c_enable_132), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n6614));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_2799.GSR = "ENABLED";
    LUT4 LM32D_CTI_O_0__bdd_1_lut (.A(dcache_refill_request), .Z(n38964)) /* synthesis lut_function=(!(A)) */ ;
    defparam LM32D_CTI_O_0__bdd_1_lut.init = 16'h5555;
    FD1P3DX creset_2795 (.D(n36326), .SP(REF_CLK_c_enable_161), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n6609));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_2795.GSR = "ENABLED";
    CCU2C add_22479_11 (.A0(adder_result_x[25]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(adder_result_x[26]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n27441), .COUT(n27442));
    defparam add_22479_11.INIT0 = 16'h5555;
    defparam add_22479_11.INIT1 = 16'h5555;
    defparam add_22479_11.INJECT1_0 = "NO";
    defparam add_22479_11.INJECT1_1 = "NO";
    FD1P3DX creset_2791 (.D(n36328), .SP(REF_CLK_c_enable_158), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n6604));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_2791.GSR = "ENABLED";
    DPR16X4C registers2 (.DI0(w_result[24]), .DI1(w_result[25]), .DI2(w_result[26]), 
            .DI3(w_result[27]), .WAD0(n45103), .WAD1(n45099), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n7610), .RAD0(n41350), 
            .RAD1(n41354), .RAD2(n41351), .RAD3(n41353), .DO0(n7569), 
            .DO1(n7570), .DO2(n7571), .DO3(n7572));
    defparam registers2.initval = "0x0000000000000000";
    FD1P3DX creset_2787 (.D(n36329), .SP(REF_CLK_c_enable_158), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n6599));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_2787.GSR = "ENABLED";
    FD1P3DX creset_2783 (.D(n36330), .SP(REF_CLK_c_enable_158), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n6594));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_2783.GSR = "ENABLED";
    FD1P3DX creset_2779 (.D(n36331), .SP(REF_CLK_c_enable_161), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n6589));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_2779.GSR = "ENABLED";
    FD1P3DX creset_2775 (.D(n36332), .SP(REF_CLK_c_enable_164), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n6584));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_2775.GSR = "ENABLED";
    FD1P3DX creset_2771 (.D(n36333), .SP(REF_CLK_c_enable_177), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n6579));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_2771.GSR = "ENABLED";
    FD1P3DX creset_2679 (.D(n36334), .SP(REF_CLK_c_enable_176), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n6434));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_2679.GSR = "ENABLED";
    FD1P3DX creset_2767 (.D(n36335), .SP(REF_CLK_c_enable_177), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n6574));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_2767.GSR = "ENABLED";
    CCU2C add_22479_15 (.A0(adder_result_x[29]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(adder_result_x[30]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n27443), .COUT(n27444));
    defparam add_22479_15.INIT0 = 16'h5555;
    defparam add_22479_15.INIT1 = 16'h5555;
    defparam add_22479_15.INJECT1_0 = "NO";
    defparam add_22479_15.INJECT1_1 = "NO";
    CCU2C add_22479_13 (.A0(adder_result_x[27]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(adder_result_x[28]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n27442), .COUT(n27443));
    defparam add_22479_13.INIT0 = 16'h5555;
    defparam add_22479_13.INIT1 = 16'h5555;
    defparam add_22479_13.INJECT1_0 = "NO";
    defparam add_22479_13.INJECT1_1 = "NO";
    LUT4 i30489_2_lut_4_lut (.A(LM32I_ADR_O[12]), .B(n45076), .C(n41390), 
         .D(SHAREDBUS_ADR_I[29]), .Z(n35647)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i30489_2_lut_4_lut.init = 16'hffca;
    LUT4 i1_2_lut_4_lut (.A(LM32I_ADR_O[12]), .B(n45076), .C(n41390), 
         .D(SHAREDBUS_ADR_I[22]), .Z(n32312)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hffca;
    LUT4 i1_2_lut_rep_858_4_lut (.A(LM32I_ADR_O[12]), .B(n45076), .C(n41390), 
         .D(SHAREDBUS_ADR_I[23]), .Z(n41263)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i1_2_lut_rep_858_4_lut.init = 16'hffca;
    DPR16X4C n66410 (.DI0(n41425), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
            .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n6637), .RAD0(n41355), 
            .RAD1(n41358), .RAD2(n41359), .RAD3(n41356), .DO0(n6642));
    defparam n66410.initval = "0x0000000000000000";
    LUT4 i1_2_lut_4_lut_adj_1043 (.A(LM32I_ADR_O[12]), .B(n45076), .C(n41390), 
         .D(n41310), .Z(n34242)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i1_2_lut_4_lut_adj_1043.init = 16'hffca;
    LUT4 i32062_3_lut (.A(n6624), .B(n6629), .C(write_idx_w[0]), .Z(n37234)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32062_3_lut.init = 16'hcaca;
    DPR16X4C n65140 (.DI0(write_idx_w[4]), .DI1(GND_net), .DI2(GND_net), 
            .DI3(GND_net), .WAD0(n45103), .WAD1(n45099), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n6640), .RAD0(n41350), 
            .RAD1(n41354), .RAD2(n41351), .RAD3(n41353), .DO0(n6515));
    defparam n65140.initval = "0x0000000000000000";
    DPR16X4C registers1 (.DI0(w_result[28]), .DI1(w_result[29]), .DI2(w_result[30]), 
            .DI3(w_result[31]), .WAD0(n45103), .WAD1(n45099), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n7610), .RAD0(n41350), 
            .RAD1(n41354), .RAD2(n41351), .RAD3(n41353), .DO0(n7573), 
            .DO1(n7574), .DO2(n7575), .DO3(n7576));
    defparam registers1.initval = "0x0000000000000000";
    LUT4 i32061_3_lut (.A(n6614), .B(n6619), .C(write_idx_w[0]), .Z(n37233)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32061_3_lut.init = 16'hcaca;
    LUT4 LM32D_CTI_O_0__bdd_4_lut (.A(LM32D_CTI_O[0]), .B(n41380), .C(locked_N_493), 
         .D(next_cycle_type_adj_6725[2]), .Z(n38963)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A (B (C (D)))) */ ;
    defparam LM32D_CTI_O_0__bdd_4_lut.init = 16'hea2a;
    LUT4 i32060_3_lut (.A(n6604), .B(n6609), .C(write_idx_w[0]), .Z(n37232)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32060_3_lut.init = 16'hcaca;
    LUT4 i32059_3_lut (.A(n6594), .B(n6599), .C(write_idx_w[0]), .Z(n37231)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32059_3_lut.init = 16'hcaca;
    DPR16X4C registers_d02 (.DI0(w_result[24]), .DI1(w_result[25]), .DI2(w_result[26]), 
            .DI3(w_result[27]), .WAD0(n45103), .WAD1(n45099), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n7610), .RAD0(n41355), 
            .RAD1(n41358), .RAD2(n41359), .RAD3(n41356), .DO0(n7637), 
            .DO1(n7638), .DO2(n7639), .DO3(n7640));
    defparam registers_d02.initval = "0x0000000000000000";
    DPR16X4C registers_d03 (.DI0(w_result[20]), .DI1(w_result[21]), .DI2(w_result[22]), 
            .DI3(w_result[23]), .WAD0(n45103), .WAD1(n45099), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n7610), .RAD0(n41355), 
            .RAD1(n41358), .RAD2(n41359), .RAD3(n41356), .DO0(n7633), 
            .DO1(n7634), .DO2(n7635), .DO3(n7636));
    defparam registers_d03.initval = "0x0000000000000000";
    DPR16X4C registers_d04 (.DI0(w_result[16]), .DI1(w_result[17]), .DI2(w_result[18]), 
            .DI3(w_result[19]), .WAD0(n45103), .WAD1(n45099), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n7610), .RAD0(n41355), 
            .RAD1(n41358), .RAD2(n41359), .RAD3(n41356), .DO0(n7629), 
            .DO1(n7630), .DO2(n7631), .DO3(n7632));
    defparam registers_d04.initval = "0x0000000000000000";
    DPR16X4C registers_d05 (.DI0(w_result[12]), .DI1(w_result[13]), .DI2(w_result[14]), 
            .DI3(w_result[15]), .WAD0(n45103), .WAD1(n45099), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n7610), .RAD0(n41355), 
            .RAD1(n41358), .RAD2(n41359), .RAD3(n41356), .DO0(n7625), 
            .DO1(n7626), .DO2(n7627), .DO3(n7628));
    defparam registers_d05.initval = "0x0000000000000000";
    DPR16X4C registers_d06 (.DI0(w_result[8]), .DI1(w_result[9]), .DI2(w_result[10]), 
            .DI3(w_result[11]), .WAD0(n45103), .WAD1(n45099), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n7610), .RAD0(n41355), 
            .RAD1(n41358), .RAD2(n41359), .RAD3(n41356), .DO0(n7621), 
            .DO1(n7622), .DO2(n7623), .DO3(n7624));
    defparam registers_d06.initval = "0x0000000000000000";
    DPR16X4C registers_d07 (.DI0(w_result[4]), .DI1(w_result[5]), .DI2(w_result[6]), 
            .DI3(w_result[7]), .WAD0(n45103), .WAD1(n45099), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n7610), .RAD0(n41355), 
            .RAD1(n41358), .RAD2(n41359), .RAD3(n41356), .DO0(n7617), 
            .DO1(n7618), .DO2(n7619), .DO3(n7620));
    defparam registers_d07.initval = "0x0000000000000000";
    DPR16X4C registers_d08 (.DI0(w_result[0]), .DI1(w_result[1]), .DI2(w_result[2]), 
            .DI3(w_result[3]), .WAD0(n45103), .WAD1(n45099), .WAD2(write_idx_w[2]), 
            .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), .WRE(n7610), .RAD0(n41355), 
            .RAD1(n41358), .RAD2(n41359), .RAD3(n41356), .DO0(n7613), 
            .DO1(n7614), .DO2(n7615), .DO3(n7616));
    defparam registers_d08.initval = "0x0000000000000000";
    DPR16X4C registers_d09 (.DI0(w_result[24]), .DI1(w_result[25]), .DI2(w_result[26]), 
            .DI3(w_result[27]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n7611), .RAD0(n41355), .RAD1(n41358), .RAD2(n41359), 
            .RAD3(n41356), .DO0(n7669), .DO1(n7670), .DO2(n7671), .DO3(n7672));
    defparam registers_d09.initval = "0x0000000000000000";
    DPR16X4C registers_d010 (.DI0(w_result[20]), .DI1(w_result[21]), .DI2(w_result[22]), 
            .DI3(w_result[23]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n7611), .RAD0(n41355), .RAD1(n41358), .RAD2(n41359), 
            .RAD3(n41356), .DO0(n7665), .DO1(n7666), .DO2(n7667), .DO3(n7668));
    defparam registers_d010.initval = "0x0000000000000000";
    DPR16X4C registers_d011 (.DI0(w_result[16]), .DI1(w_result[17]), .DI2(w_result[18]), 
            .DI3(w_result[19]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n7611), .RAD0(n41355), .RAD1(n41358), .RAD2(n41359), 
            .RAD3(n41356), .DO0(n7661), .DO1(n7662), .DO2(n7663), .DO3(n7664));
    defparam registers_d011.initval = "0x0000000000000000";
    DPR16X4C registers_d012 (.DI0(w_result[12]), .DI1(w_result[13]), .DI2(w_result[14]), 
            .DI3(w_result[15]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n7611), .RAD0(n41355), .RAD1(n41358), .RAD2(n41359), 
            .RAD3(n41356), .DO0(n7657), .DO1(n7658), .DO2(n7659), .DO3(n7660));
    defparam registers_d012.initval = "0x0000000000000000";
    DPR16X4C registers_d013 (.DI0(w_result[8]), .DI1(w_result[9]), .DI2(w_result[10]), 
            .DI3(w_result[11]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n7611), .RAD0(n41355), .RAD1(n41358), .RAD2(n41359), 
            .RAD3(n41356), .DO0(n7653), .DO1(n7654), .DO2(n7655), .DO3(n7656));
    defparam registers_d013.initval = "0x0000000000000000";
    DPR16X4C registers_d014 (.DI0(w_result[4]), .DI1(w_result[5]), .DI2(w_result[6]), 
            .DI3(w_result[7]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n7611), .RAD0(n41355), .RAD1(n41358), .RAD2(n41359), 
            .RAD3(n41356), .DO0(n7649), .DO1(n7650), .DO2(n7651), .DO3(n7652));
    defparam registers_d014.initval = "0x0000000000000000";
    DPR16X4C registers_d015 (.DI0(w_result[0]), .DI1(w_result[1]), .DI2(w_result[2]), 
            .DI3(w_result[3]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(REF_CLK_c), 
            .WRE(n7611), .RAD0(n41355), .RAD1(n41358), .RAD2(n41359), 
            .RAD3(n41356), .DO0(n7645), .DO1(n7646), .DO2(n7647), .DO3(n7648));
    defparam registers_d015.initval = "0x0000000000000000";
    IB USER_BUTTON_pad (.I(USER_BUTTON), .O(USER_BUTTON_c));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(24[7:18])
    IB REF_CLK_pad (.I(REF_CLK), .O(REF_CLK_c));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    OB IO_0_pad (.I(IO_0_c_0), .O(IO_0));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(31[3:7])
    OB IO_MISO_pad (.I(IO_MISO_c), .O(IO_MISO));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(30[3:10])
    OB IO_MOSI_pad (.I(IO_MOSI_c), .O(IO_MOSI));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(29[3:10])
    OB IO_SCK_pad (.I(IO_SCK_c), .O(IO_SCK));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(28[3:9])
    OB LED_B_pad (.I(LED_B_c_0), .O(LED_B));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(27[3:8])
    OB LED_G_pad (.I(LED_G_c_0), .O(LED_G));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(26[3:8])
    OB LED_R_pad (.I(LED_R_c_0), .O(LED_R));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(25[7:12])
    LUT4 i32058_3_lut (.A(n6584), .B(n6589), .C(write_idx_w[0]), .Z(n37230)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32058_3_lut.init = 16'hcaca;
    LUT4 i32057_3_lut (.A(n6574), .B(n6579), .C(write_idx_w[0]), .Z(n37229)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32057_3_lut.init = 16'hcaca;
    LUT4 i32056_3_lut (.A(n6434), .B(n6439), .C(write_idx_w[0]), .Z(n37228)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32056_3_lut.init = 16'hcaca;
    CCU2C add_22479_5 (.A0(adder_result_x[19]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(adder_result_x[20]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n27438), .COUT(n27439));
    defparam add_22479_5.INIT0 = 16'h5555;
    defparam add_22479_5.INIT1 = 16'h5555;
    defparam add_22479_5.INJECT1_0 = "NO";
    defparam add_22479_5.INJECT1_1 = "NO";
    LUT4 i32055_3_lut (.A(n6424), .B(n6429), .C(write_idx_w[0]), .Z(n37227)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32055_3_lut.init = 16'hcaca;
    CCU2C add_22479_3 (.A0(adder_result_x[17]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(adder_result_x[18]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n27437), .COUT(n27438));
    defparam add_22479_3.INIT0 = 16'h5555;
    defparam add_22479_3.INIT1 = 16'h5555;
    defparam add_22479_3.INJECT1_0 = "NO";
    defparam add_22479_3.INJECT1_1 = "NO";
    PFUMX i32337 (.BLUT(n37507), .ALUT(n37508), .C0(n41356), .Z(n37509));
    PFUMX i32012 (.BLUT(n37176), .ALUT(n37177), .C0(n41354), .Z(n37184));
    PFUMX i32013 (.BLUT(n37178), .ALUT(n37179), .C0(n41354), .Z(n37185));
    PFUMX i32014 (.BLUT(n37180), .ALUT(n37181), .C0(n41354), .Z(n37186));
    PFUMX i32015 (.BLUT(n37182), .ALUT(n37183), .C0(n41354), .Z(n37187));
    PFUMX i32069 (.BLUT(n37239), .ALUT(n37240), .C0(write_idx_w[3]), .Z(n6502));
    PFUMX i32331 (.BLUT(n37495), .ALUT(n37496), .C0(n41358), .Z(n37503));
    PFUMX i32332 (.BLUT(n37497), .ALUT(n37498), .C0(n41358), .Z(n37504));
    PFUMX i32333 (.BLUT(n37499), .ALUT(n37500), .C0(n41358), .Z(n37505));
    PFUMX i32334 (.BLUT(n37501), .ALUT(n37502), .C0(n41358), .Z(n37506));
    CCU2C _add_1_3756_add_4_9 (.A0(flush_set[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(flush_set[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n27508), .S0(flush_set_8__N_1953[7]), .S1(flush_set_8__N_1953[8]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(421[29:45])
    defparam _add_1_3756_add_4_9.INIT0 = 16'h555f;
    defparam _add_1_3756_add_4_9.INIT1 = 16'h555f;
    defparam _add_1_3756_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3756_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3756_add_4_7 (.A0(flush_set[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(flush_set[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n27507), .COUT(n27508), .S0(flush_set_8__N_1953[5]), 
          .S1(flush_set_8__N_1953[6]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(421[29:45])
    defparam _add_1_3756_add_4_7.INIT0 = 16'h555f;
    defparam _add_1_3756_add_4_7.INIT1 = 16'h555f;
    defparam _add_1_3756_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3756_add_4_7.INJECT1_1 = "NO";
    LUT4 i1_3_lut (.A(write_idx_w[1]), .B(n41325), .C(write_idx_w[0]), 
         .Z(REF_CLK_c_enable_161)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    CCU2C _add_1_3756_add_4_5 (.A0(flush_set[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(flush_set[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n27506), .COUT(n27507), .S0(flush_set_8__N_1953[3]), 
          .S1(flush_set_8__N_1953[4]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(421[29:45])
    defparam _add_1_3756_add_4_5.INIT0 = 16'h555f;
    defparam _add_1_3756_add_4_5.INIT1 = 16'h555f;
    defparam _add_1_3756_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3756_add_4_5.INJECT1_1 = "NO";
    PFUMX i34383 (.BLUT(n41495), .ALUT(n41496), .C0(n45101), .Z(n29));
    CCU2C _add_1_3756_add_4_3 (.A0(flush_set[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(flush_set[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n27505), .COUT(n27506), .S0(flush_set_8__N_1953[1]), 
          .S1(flush_set_8__N_1953[2]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(421[29:45])
    defparam _add_1_3756_add_4_3.INIT0 = 16'h555f;
    defparam _add_1_3756_add_4_3.INIT1 = 16'h555f;
    defparam _add_1_3756_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3756_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3756_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(flush_set[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n27505), .S1(flush_set_8__N_1953[0]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(421[29:45])
    defparam _add_1_3756_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3756_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3756_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3756_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_9 (.A0(flush_set_adj_6801[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(flush_set_adj_6801[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n27503), .S0(flush_set_8__N_2513[7]), 
          .S1(flush_set_8__N_2513[8]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(483[29:45])
    defparam _add_1_3753_add_4_9.INIT0 = 16'h555f;
    defparam _add_1_3753_add_4_9.INIT1 = 16'h555f;
    defparam _add_1_3753_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_7 (.A0(flush_set_adj_6801[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(flush_set_adj_6801[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n27502), .COUT(n27503), .S0(flush_set_8__N_2513[5]), 
          .S1(flush_set_8__N_2513[6]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(483[29:45])
    defparam _add_1_3753_add_4_7.INIT0 = 16'h555f;
    defparam _add_1_3753_add_4_7.INIT1 = 16'h555f;
    defparam _add_1_3753_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_5 (.A0(flush_set_adj_6801[3]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(flush_set_adj_6801[4]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n27501), .COUT(n27502), .S0(flush_set_8__N_2513[3]), 
          .S1(flush_set_8__N_2513[4]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(483[29:45])
    defparam _add_1_3753_add_4_5.INIT0 = 16'h555f;
    defparam _add_1_3753_add_4_5.INIT1 = 16'h555f;
    defparam _add_1_3753_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3753_add_4_3 (.A0(flush_set_adj_6801[1]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(flush_set_adj_6801[2]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n27500), .COUT(n27501), .S0(flush_set_8__N_2513[1]), 
          .S1(flush_set_8__N_2513[2]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(483[29:45])
    defparam _add_1_3753_add_4_3.INIT0 = 16'h555f;
    defparam _add_1_3753_add_4_3.INIT1 = 16'h555f;
    defparam _add_1_3753_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_3.INJECT1_1 = "NO";
    LUT4 i31164_4_lut (.A(dc_re), .B(operand_1_x[1]), .C(n41379), .D(n41394), 
         .Z(n36336)) /* synthesis lut_function=(A (B+(C+(D)))+!A !((C+(D))+!B)) */ ;
    defparam i31164_4_lut.init = 16'haaac;
    CCU2C _add_1_3753_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(flush_set_adj_6801[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n27500), .S1(flush_set_8__N_2513[0]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(483[29:45])
    defparam _add_1_3753_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3753_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3753_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3753_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_31 (.A0(pc_d[31]), .B0(n6781), .C0(n45106), 
          .D0(n34), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27499), .S0(branch_target_d[31]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam _add_1_3750_add_4_31.INIT0 = 16'h9aaa;
    defparam _add_1_3750_add_4_31.INIT1 = 16'h0000;
    defparam _add_1_3750_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_31.INJECT1_1 = "NO";
    LUT4 i8_3_lut (.A(\genblk1.pmi_address [12]), .B(n41303), .C(n20000), 
         .Z(\genblk1.read_address [10])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i8_3_lut.init = 16'hacac;
    LUT4 i12_3_lut (.A(n41303), .B(\genblk1.pmi_address [12]), .C(n6038), 
         .Z(\genblk1.write_address [10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12_3_lut.init = 16'hcaca;
    CCU2C _add_1_3750_add_4_29 (.A0(pc_d[29]), .B0(n6781), .C0(n45106), 
          .D0(n34), .A1(pc_d[30]), .B1(n6781), .C1(n45106), .D1(n34), 
          .CIN(n27498), .COUT(n27499), .S0(branch_target_d[29]), .S1(branch_target_d[30]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam _add_1_3750_add_4_29.INIT0 = 16'h9aaa;
    defparam _add_1_3750_add_4_29.INIT1 = 16'h9aaa;
    defparam _add_1_3750_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_27 (.A0(pc_d[27]), .B0(n6781), .C0(n45105), 
          .D0(n34), .A1(pc_d[28]), .B1(n6781), .C1(n45105), .D1(n34), 
          .CIN(n27497), .COUT(n27498), .S0(branch_target_d[27]), .S1(branch_target_d[28]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam _add_1_3750_add_4_27.INIT0 = 16'h9aaa;
    defparam _add_1_3750_add_4_27.INIT1 = 16'h9aaa;
    defparam _add_1_3750_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_27.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_25 (.A0(pc_d[25]), .B0(n6781), .C0(n45106), 
          .D0(n36), .A1(pc_d[26]), .B1(n6781), .C1(n45106), .D1(n37), 
          .CIN(n27496), .COUT(n27497), .S0(branch_target_d[25]), .S1(branch_target_d[26]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam _add_1_3750_add_4_25.INIT0 = 16'h9aaa;
    defparam _add_1_3750_add_4_25.INIT1 = 16'h9aaa;
    defparam _add_1_3750_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_23 (.A0(pc_d[23]), .B0(n6781), .C0(n10593), 
          .D0(n45106), .A1(pc_d[24]), .B1(n6781), .C1(n10595), .D1(n45106), 
          .CIN(n27495), .COUT(n27496), .S0(branch_target_d[23]), .S1(branch_target_d[24]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam _add_1_3750_add_4_23.INIT0 = 16'h9aaa;
    defparam _add_1_3750_add_4_23.INIT1 = 16'h9aaa;
    defparam _add_1_3750_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_21 (.A0(pc_d[21]), .B0(n6781), .C0(n10589), 
          .D0(n45106), .A1(pc_d[22]), .B1(n6781), .C1(n10591), .D1(n45106), 
          .CIN(n27494), .COUT(n27495), .S0(branch_target_d[21]), .S1(branch_target_d[22]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam _add_1_3750_add_4_21.INIT0 = 16'h9aaa;
    defparam _add_1_3750_add_4_21.INIT1 = 16'h9aaa;
    defparam _add_1_3750_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_19 (.A0(pc_d[19]), .B0(n6781), .C0(n10585), 
          .D0(n45106), .A1(pc_d[20]), .B1(n6781), .C1(n10587), .D1(n45106), 
          .CIN(n27493), .COUT(n27494), .S0(branch_target_d[19]), .S1(branch_target_d[20]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam _add_1_3750_add_4_19.INIT0 = 16'h9aaa;
    defparam _add_1_3750_add_4_19.INIT1 = 16'h9aaa;
    defparam _add_1_3750_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_17 (.A0(pc_d[17]), .B0(n6781), .C0(n6764), 
          .D0(n45106), .A1(pc_d[18]), .B1(n6781), .C1(n10452), .D1(n45106), 
          .CIN(n27492), .COUT(n27493), .S0(branch_target_d[17]), .S1(branch_target_d[18]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam _add_1_3750_add_4_17.INIT0 = 16'h9aaa;
    defparam _add_1_3750_add_4_17.INIT1 = 16'h9aaa;
    defparam _add_1_3750_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_15 (.A0(pc_d[15]), .B0(n6781), .C0(n45106), 
          .D0(n6762), .A1(pc_d[16]), .B1(n6781), .C1(n45106), .D1(n6763), 
          .CIN(n27491), .COUT(n27492), .S0(branch_target_d[15]), .S1(branch_target_d[16]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam _add_1_3750_add_4_15.INIT0 = 16'h9aaa;
    defparam _add_1_3750_add_4_15.INIT1 = 16'h9aaa;
    defparam _add_1_3750_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_13 (.A0(pc_d[13]), .B0(n6781), .C0(n45106), 
          .D0(n6760), .A1(pc_d[14]), .B1(n6781), .C1(n45106), .D1(n6761), 
          .CIN(n27490), .COUT(n27491), .S0(branch_target_d[13]), .S1(branch_target_d[14]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam _add_1_3750_add_4_13.INIT0 = 16'h9aaa;
    defparam _add_1_3750_add_4_13.INIT1 = 16'h9aaa;
    defparam _add_1_3750_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_11 (.A0(pc_d[11]), .B0(n6781), .C0(n6758), 
          .D0(n45106), .A1(pc_d[12]), .B1(n6781), .C1(n6759), .D1(n45106), 
          .CIN(n27489), .COUT(n27490), .S0(branch_target_d[11]), .S1(branch_target_d[12]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam _add_1_3750_add_4_11.INIT0 = 16'h9aaa;
    defparam _add_1_3750_add_4_11.INIT1 = 16'h9aaa;
    defparam _add_1_3750_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_11.INJECT1_1 = "NO";
    LUT4 i2815_3_lut (.A(write_idx_w[4]), .B(n41325), .C(n6502), .Z(n6637)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i2815_3_lut.init = 16'h4c4c;
    LUT4 i2818_3_lut (.A(write_idx_w[4]), .B(n41325), .C(n6502), .Z(n6640)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i2818_3_lut.init = 16'h8c8c;
    CCU2C _add_1_3750_add_4_9 (.A0(pc_d[9]), .B0(n6781), .C0(n6756), .D0(n45106), 
          .A1(pc_d[10]), .B1(n6781), .C1(n6757), .D1(n45106), .CIN(n27488), 
          .COUT(n27489), .S0(branch_target_d[9]), .S1(branch_target_d[10]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam _add_1_3750_add_4_9.INIT0 = 16'h9aaa;
    defparam _add_1_3750_add_4_9.INIT1 = 16'h9aaa;
    defparam _add_1_3750_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_7 (.A0(pc_d[7]), .B0(n6781), .C0(n6754), .D0(n45106), 
          .A1(pc_d[8]), .B1(n6781), .C1(n6755), .D1(n45106), .CIN(n27487), 
          .COUT(n27488), .S0(branch_target_d[7]), .S1(branch_target_d[8]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam _add_1_3750_add_4_7.INIT0 = 16'h9aaa;
    defparam _add_1_3750_add_4_7.INIT1 = 16'h9aaa;
    defparam _add_1_3750_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_5 (.A0(pc_d[5]), .B0(n6781), .C0(n6752), .D0(n45106), 
          .A1(pc_d[6]), .B1(n6781), .C1(n6753), .D1(n45106), .CIN(n27486), 
          .COUT(n27487), .S0(branch_target_d[5]), .S1(branch_target_d[6]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam _add_1_3750_add_4_5.INIT0 = 16'h9aaa;
    defparam _add_1_3750_add_4_5.INIT1 = 16'h9aaa;
    defparam _add_1_3750_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_3 (.A0(pc_d[3]), .B0(n6781), .C0(n6750), .D0(n45106), 
          .A1(pc_d[4]), .B1(n6781), .C1(n6751), .D1(n45106), .CIN(n27485), 
          .COUT(n27486), .S0(branch_target_d[3]), .S1(branch_target_d[4]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam _add_1_3750_add_4_3.INIT0 = 16'h9aaa;
    defparam _add_1_3750_add_4_3.INIT1 = 16'h9aaa;
    defparam _add_1_3750_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3750_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc_d[2]), .B1(n6781), .C1(n6749), .D1(n45106), 
          .COUT(n27485), .S1(branch_target_d[2]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam _add_1_3750_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3750_add_4_1.INIT1 = 16'h9aaa;
    defparam _add_1_3750_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3750_add_4_1.INJECT1_1 = "NO";
    LUT4 i12515_3_lut (.A(operand_m[5]), .B(dcache_refill_address[5]), .C(state_adj_6798[2]), 
         .Z(dmem_write_address_adj_6796[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(186[26:31])
    defparam i12515_3_lut.init = 16'hcaca;
    LUT4 i12512_3_lut (.A(operand_m[9]), .B(dcache_refill_address[9]), .C(state_adj_6798[2]), 
         .Z(dmem_write_address_adj_6796[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(186[26:31])
    defparam i12512_3_lut.init = 16'hcaca;
    LUT4 i12511_3_lut (.A(operand_m[10]), .B(dcache_refill_address[10]), 
         .C(state_adj_6798[2]), .Z(dmem_write_address_adj_6796[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(186[26:31])
    defparam i12511_3_lut.init = 16'hcaca;
    LUT4 i12514_3_lut (.A(dcache_refill_address[5]), .B(flush_set_adj_6801[1]), 
         .C(state_adj_6798[0]), .Z(tmem_write_address_adj_6794[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(186[26:31])
    defparam i12514_3_lut.init = 16'hcaca;
    LUT4 i31165_4_lut (.A(bie), .B(bie_N_3274), .C(n31279), .D(n41401), 
         .Z(n36337)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;
    defparam i31165_4_lut.init = 16'hccca;
    CCU2C _add_1_3765_add_4_15 (.A0(n11843), .B0(\genblk1.state [2]), .C0(\genblk1.pmi_address [13]), 
          .D0(n41300), .A1(n11843), .B1(\genblk1.state [2]), .C1(\genblk1.pmi_address [14]), 
          .D1(n41298), .CIN(n27483), .S0(n37_adj_6598), .S1(n34_adj_6597));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(434[7] 442[10])
    defparam _add_1_3765_add_4_15.INIT0 = 16'hf1e0;
    defparam _add_1_3765_add_4_15.INIT1 = 16'hf1e0;
    defparam _add_1_3765_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_15.INJECT1_1 = "NO";
    LUT4 i12518_3_lut (.A(dcache_refill_address[9]), .B(flush_set_adj_6801[5]), 
         .C(state_adj_6798[0]), .Z(tmem_write_address_adj_6794[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(186[26:31])
    defparam i12518_3_lut.init = 16'hcaca;
    CCU2C _add_1_3765_add_4_13 (.A0(n11843), .B0(\genblk1.state [2]), .C0(\genblk1.pmi_address [11]), 
          .D0(n41299), .A1(n11843), .B1(\genblk1.state [2]), .C1(\genblk1.pmi_address [12]), 
          .D1(n41303), .CIN(n27482), .COUT(n27483), .S0(n43), .S1(n40));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(434[7] 442[10])
    defparam _add_1_3765_add_4_13.INIT0 = 16'hf1e0;
    defparam _add_1_3765_add_4_13.INIT1 = 16'hf1e0;
    defparam _add_1_3765_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_13.INJECT1_1 = "NO";
    LUT4 i12517_3_lut (.A(dcache_refill_address[10]), .B(flush_set_adj_6801[6]), 
         .C(state_adj_6798[0]), .Z(tmem_write_address_adj_6794[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(186[26:31])
    defparam i12517_3_lut.init = 16'hcaca;
    CCU2C _add_1_3765_add_4_11 (.A0(n11843), .B0(\genblk1.state [2]), .C0(\genblk1.pmi_address [9]), 
          .D0(n41310), .A1(n11843), .B1(\genblk1.state [2]), .C1(\genblk1.pmi_address [10]), 
          .D1(SHAREDBUS_ADR_I[10]), .CIN(n27481), .COUT(n27482), .S0(n49), 
          .S1(n46));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(434[7] 442[10])
    defparam _add_1_3765_add_4_11.INIT0 = 16'hf1e0;
    defparam _add_1_3765_add_4_11.INIT1 = 16'hf1e0;
    defparam _add_1_3765_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_9 (.A0(n11843), .B0(\genblk1.state [2]), .C0(\genblk1.pmi_address [7]), 
          .D0(SHAREDBUS_ADR_I[7]), .A1(n11843), .B1(\genblk1.state [2]), 
          .C1(\genblk1.pmi_address [8]), .D1(n41301), .CIN(n27480), .COUT(n27481), 
          .S0(n55), .S1(n52));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(434[7] 442[10])
    defparam _add_1_3765_add_4_9.INIT0 = 16'hf1e0;
    defparam _add_1_3765_add_4_9.INIT1 = 16'hf1e0;
    defparam _add_1_3765_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_7 (.A0(n11843), .B0(\genblk1.state [2]), .C0(\genblk1.pmi_address [5]), 
          .D0(SHAREDBUS_ADR_I[5]), .A1(n11843), .B1(\genblk1.state [2]), 
          .C1(\genblk1.pmi_address [6]), .D1(n41346), .CIN(n27479), .COUT(n27480), 
          .S0(n61), .S1(n58));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(434[7] 442[10])
    defparam _add_1_3765_add_4_7.INIT0 = 16'hf1e0;
    defparam _add_1_3765_add_4_7.INIT1 = 16'hf1e0;
    defparam _add_1_3765_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_5 (.A0(n11843), .B0(\genblk1.state [2]), .C0(\genblk1.pmi_address [3]), 
          .D0(n41344), .A1(n11843), .B1(\genblk1.state [2]), .C1(\genblk1.pmi_address [4]), 
          .D1(n41347), .CIN(n27478), .COUT(n27479), .S0(n67_adj_6600), 
          .S1(n64_adj_6599));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(434[7] 442[10])
    defparam _add_1_3765_add_4_5.INIT0 = 16'hf1e0;
    defparam _add_1_3765_add_4_5.INIT1 = 16'hf1e0;
    defparam _add_1_3765_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_3 (.A0(n3485), .B0(n5386), .C0(n3700), .D0(n41321), 
          .A1(n3432), .B1(n6034), .C1(n41292), .D1(n19822), .CIN(n27477), 
          .COUT(n27478), .S0(n73_adj_6602), .S1(n70_adj_6601));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(434[7] 442[10])
    defparam _add_1_3765_add_4_3.INIT0 = 16'h2112;
    defparam _add_1_3765_add_4_3.INIT1 = 16'h9aaa;
    defparam _add_1_3765_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3765_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n5085), .B1(n6034), .C1(n8), .D1(n3486), 
          .COUT(n27477), .S1(n76_adj_6603));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(434[7] 442[10])
    defparam _add_1_3765_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3765_add_4_1.INIT1 = 16'h65aa;
    defparam _add_1_3765_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3765_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_31 (.A0(pc_f[31]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27476), .S0(n64));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[13:24])
    defparam _add_1_3759_add_4_31.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_31.INIT1 = 16'h0000;
    defparam _add_1_3759_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_29 (.A0(pc_f[29]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc_f[30]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n27475), .COUT(n27476), .S0(n70), .S1(n67));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[13:24])
    defparam _add_1_3759_add_4_29.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_29.INIT1 = 16'haaa0;
    defparam _add_1_3759_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_27 (.A0(pc_f[27]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc_f[28]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n27474), .COUT(n27475), .S0(n76), .S1(n73));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[13:24])
    defparam _add_1_3759_add_4_27.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_27.INIT1 = 16'haaa0;
    defparam _add_1_3759_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_27.INJECT1_1 = "NO";
    LUT4 i33427_then_3_lut (.A(LM32D_ADR_O[19]), .B(selected[0]), .C(LM32D_ADR_O[17]), 
         .Z(n41496)) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;
    defparam i33427_then_3_lut.init = 16'h3232;
    LUT4 i33427_else_3_lut (.A(LM32I_ADR_O[17]), .B(LM32I_ADR_O[19]), .C(selected[0]), 
         .Z(n41495)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i33427_else_3_lut.init = 16'he0e0;
    LUT4 i12513_3_lut (.A(operand_m[5]), .B(dcache_refill_address[5]), .C(dcache_refill_request), 
         .Z(d_adr_o_31__N_2278[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(676[6:27])
    defparam i12513_3_lut.init = 16'hcaca;
    LUT4 i12516_3_lut (.A(operand_m[9]), .B(dcache_refill_address[9]), .C(dcache_refill_request), 
         .Z(d_adr_o_31__N_2278[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(676[6:27])
    defparam i12516_3_lut.init = 16'hcaca;
    LUT4 i12510_3_lut (.A(operand_m[10]), .B(dcache_refill_address[10]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(676[6:27])
    defparam i12510_3_lut.init = 16'hcaca;
    CCU2C _add_1_3759_add_4_25 (.A0(pc_f[25]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc_f[26]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n27473), .COUT(n27474), .S0(n82), .S1(n79));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[13:24])
    defparam _add_1_3759_add_4_25.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_25.INIT1 = 16'haaa0;
    defparam _add_1_3759_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_23 (.A0(pc_f[23]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc_f[24]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n27472), .COUT(n27473), .S0(n88), .S1(n85));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[13:24])
    defparam _add_1_3759_add_4_23.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_23.INIT1 = 16'haaa0;
    defparam _add_1_3759_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_21 (.A0(pc_f[21]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc_f[22]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n27471), .COUT(n27472), .S0(n94), .S1(n91));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[13:24])
    defparam _add_1_3759_add_4_21.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_21.INIT1 = 16'haaa0;
    defparam _add_1_3759_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_19 (.A0(pc_f[19]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc_f[20]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n27470), .COUT(n27471), .S0(n100), .S1(n97));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[13:24])
    defparam _add_1_3759_add_4_19.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_3759_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_17 (.A0(pc_f[17]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc_f[18]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n27469), .COUT(n27470), .S0(n106), .S1(n103));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[13:24])
    defparam _add_1_3759_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_17.INIT1 = 16'haaa0;
    defparam _add_1_3759_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_17.INJECT1_1 = "NO";
    LUT4 i33099_2_lut_rep_990 (.A(write_idx_w[2]), .B(write_idx_w[3]), .Z(REF_CLK_c_enable_177)) /* synthesis lut_function=(!((B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i33099_2_lut_rep_990.init = 16'h2222;
    LUT4 i31160_3_lut_3_lut (.A(write_idx_w[2]), .B(write_idx_w[3]), .C(n6584), 
         .Z(n36332)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i31160_3_lut_3_lut.init = 16'hf2f2;
    LUT4 i31159_3_lut_3_lut (.A(write_idx_w[2]), .B(write_idx_w[3]), .C(n6589), 
         .Z(n36331)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i31159_3_lut_3_lut.init = 16'hf2f2;
    CCU2C _add_1_3759_add_4_15 (.A0(pc_f[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc_f[16]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n27468), .COUT(n27469), .S0(n112), .S1(n109));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[13:24])
    defparam _add_1_3759_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_3759_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_15.INJECT1_1 = "NO";
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    CCU2C _add_1_3759_add_4_13 (.A0(pc_f[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc_f[14]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n27467), .COUT(n27468), .S0(n118), .S1(n115));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[13:24])
    defparam _add_1_3759_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_3759_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_11 (.A0(pc_f[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc_f[12]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n27466), .COUT(n27467), .S0(n124), .S1(n121));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[13:24])
    defparam _add_1_3759_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_3759_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_9 (.A0(pc_f[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc_f[10]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n27465), .COUT(n27466), .S0(n130), .S1(n127));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[13:24])
    defparam _add_1_3759_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_3759_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_9.INJECT1_1 = "NO";
    PFUMX i32063 (.BLUT(n37227), .ALUT(n37228), .C0(write_idx_w[1]), .Z(n37235));
    CCU2C _add_1_3759_add_4_7 (.A0(pc_f[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc_f[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n27464), .COUT(n27465), .S0(n136), .S1(n133));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[13:24])
    defparam _add_1_3759_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_3759_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_5 (.A0(pc_f[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc_f[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n27463), .COUT(n27464), .S0(n142), .S1(n139));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[13:24])
    defparam _add_1_3759_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_3759_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_3 (.A0(pc_f[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc_f[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n27462), .COUT(n27463), .S0(n148), .S1(n145));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[13:24])
    defparam _add_1_3759_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_3759_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_3759_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_3759_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pc_f[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n27462), .S1(n151));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[13:24])
    defparam _add_1_3759_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_3759_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_3759_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_3759_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_34 (.A0(b[31]), .B0(p[30]), .C0(GND_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n27460), 
          .S0(t[31]), .S1(t[32]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam _add_1_add_4_34.INIT0 = 16'h9995;
    defparam _add_1_add_4_34.INIT1 = 16'hffff;
    defparam _add_1_add_4_34.INJECT1_0 = "NO";
    defparam _add_1_add_4_34.INJECT1_1 = "NO";
    LUT4 i990_4_lut (.A(n35448), .B(n45179), .C(IO_0_c_0), .D(n2023), 
         .Z(REF_CLK_c_enable_1424)) /* synthesis lut_function=(A (B)+!A !((C+!(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(115[7] 124[14])
    defparam i990_4_lut.init = 16'h8c88;
    CCU2C _add_1_add_4_32 (.A0(b[29]), .B0(p[28]), .C0(GND_net), .D0(VCC_net), 
          .A1(b[30]), .B1(p[29]), .C1(GND_net), .D1(VCC_net), .CIN(n27459), 
          .COUT(n27460), .S0(t[29]), .S1(t[30]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam _add_1_add_4_32.INIT0 = 16'h9995;
    defparam _add_1_add_4_32.INIT1 = 16'h9995;
    defparam _add_1_add_4_32.INJECT1_0 = "NO";
    defparam _add_1_add_4_32.INJECT1_1 = "NO";
    PFUMX i32064 (.BLUT(n37229), .ALUT(n37230), .C0(write_idx_w[1]), .Z(n37236));
    PFUMX i32065 (.BLUT(n37231), .ALUT(n37232), .C0(write_idx_w[1]), .Z(n37237));
    PFUMX i32066 (.BLUT(n37233), .ALUT(n37234), .C0(write_idx_w[1]), .Z(n37238));
    CCU2C _add_1_add_4_30 (.A0(b[27]), .B0(p[26]), .C0(GND_net), .D0(VCC_net), 
          .A1(b[28]), .B1(p[27]), .C1(GND_net), .D1(VCC_net), .CIN(n27458), 
          .COUT(n27459), .S0(t[27]), .S1(t[28]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam _add_1_add_4_30.INIT0 = 16'h9995;
    defparam _add_1_add_4_30.INIT1 = 16'h9995;
    defparam _add_1_add_4_30.INJECT1_0 = "NO";
    defparam _add_1_add_4_30.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_28 (.A0(b[25]), .B0(p[24]), .C0(GND_net), .D0(VCC_net), 
          .A1(b[26]), .B1(p[25]), .C1(GND_net), .D1(VCC_net), .CIN(n27457), 
          .COUT(n27458), .S0(t[25]), .S1(t[26]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam _add_1_add_4_28.INIT0 = 16'h9995;
    defparam _add_1_add_4_28.INIT1 = 16'h9995;
    defparam _add_1_add_4_28.INJECT1_0 = "NO";
    defparam _add_1_add_4_28.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_26 (.A0(b[23]), .B0(p[22]), .C0(GND_net), .D0(VCC_net), 
          .A1(b[24]), .B1(p[23]), .C1(GND_net), .D1(VCC_net), .CIN(n27456), 
          .COUT(n27457), .S0(t[23]), .S1(t[24]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam _add_1_add_4_26.INIT0 = 16'h9995;
    defparam _add_1_add_4_26.INIT1 = 16'h9995;
    defparam _add_1_add_4_26.INJECT1_0 = "NO";
    defparam _add_1_add_4_26.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_24 (.A0(b[21]), .B0(p[20]), .C0(GND_net), .D0(VCC_net), 
          .A1(b[22]), .B1(p[21]), .C1(GND_net), .D1(VCC_net), .CIN(n27455), 
          .COUT(n27456), .S0(t[21]), .S1(t[22]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam _add_1_add_4_24.INIT0 = 16'h9995;
    defparam _add_1_add_4_24.INIT1 = 16'h9995;
    defparam _add_1_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_22 (.A0(b[19]), .B0(p[18]), .C0(GND_net), .D0(VCC_net), 
          .A1(b[20]), .B1(p[19]), .C1(GND_net), .D1(VCC_net), .CIN(n27454), 
          .COUT(n27455), .S0(t[19]), .S1(t[20]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam _add_1_add_4_22.INIT0 = 16'h9995;
    defparam _add_1_add_4_22.INIT1 = 16'h9995;
    defparam _add_1_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_add_4_22.INJECT1_1 = "NO";
    LUT4 i15228_3_lut (.A(counter[2]), .B(n2), .C(n3), .Z(n12428)) /* synthesis lut_function=(A+(B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(472[15:29])
    defparam i15228_3_lut.init = 16'heaea;
    LUT4 i33090_2_lut_rep_998 (.A(write_idx_w[2]), .B(write_idx_w[3]), .Z(REF_CLK_c_enable_158)) /* synthesis lut_function=(!(A+!(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i33090_2_lut_rep_998.init = 16'h4444;
    LUT4 i31154_3_lut_3_lut (.A(write_idx_w[2]), .B(write_idx_w[3]), .C(n6609), 
         .Z(n36326)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i31154_3_lut_3_lut.init = 16'hf4f4;
    LUT4 equal_2673_i5_2_lut_rep_1000 (.A(write_idx_w[0]), .B(write_idx_w[1]), 
         .Z(n41405)) /* synthesis lut_function=(A+!(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam equal_2673_i5_2_lut_rep_1000.init = 16'hbbbb;
    LUT4 i31156_3_lut_3_lut_4_lut (.A(write_idx_w[0]), .B(write_idx_w[1]), 
         .C(n6604), .D(n41325), .Z(n36328)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i31156_3_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 i31162_3_lut_3_lut (.A(write_idx_w[0]), .B(write_idx_w[1]), .C(n6434), 
         .Z(n36334)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i31162_3_lut_3_lut.init = 16'hf4f4;
    LUT4 i31151_3_lut_3_lut_4_lut (.A(write_idx_w[0]), .B(write_idx_w[1]), 
         .C(n6624), .D(n41325), .Z(n36323)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i31151_3_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 i14753_2_lut_rep_1002 (.A(write_idx_w[2]), .B(write_idx_w[3]), 
         .Z(REF_CLK_c_enable_132)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14753_2_lut_rep_1002.init = 16'h8888;
    LUT4 i31150_3_lut_3_lut (.A(write_idx_w[2]), .B(write_idx_w[3]), .C(n6629), 
         .Z(n36322)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i31150_3_lut_3_lut.init = 16'hf8f8;
    CCU2C _add_1_add_4_20 (.A0(b[17]), .B0(p[16]), .C0(GND_net), .D0(VCC_net), 
          .A1(b[18]), .B1(p[17]), .C1(GND_net), .D1(VCC_net), .CIN(n27453), 
          .COUT(n27454), .S0(t[17]), .S1(t[18]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam _add_1_add_4_20.INIT0 = 16'h9995;
    defparam _add_1_add_4_20.INIT1 = 16'h9995;
    defparam _add_1_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_add_4_20.INJECT1_1 = "NO";
    LUT4 i31166_4_lut (.A(LED_R_c_0), .B(SHAREDBUS_DAT_I[24]), .C(n29830), 
         .D(n35006), .Z(n36338)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i31166_4_lut.init = 16'hcaaa;
    CCU2C _add_1_add_4_18 (.A0(b[15]), .B0(p[14]), .C0(GND_net), .D0(VCC_net), 
          .A1(b[16]), .B1(p[15]), .C1(GND_net), .D1(VCC_net), .CIN(n27452), 
          .COUT(n27453), .S0(t[15]), .S1(t[16]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam _add_1_add_4_18.INIT0 = 16'h9995;
    defparam _add_1_add_4_18.INIT1 = 16'h9995;
    defparam _add_1_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_add_4_18.INJECT1_1 = "NO";
    LUT4 i31167_4_lut (.A(LED_B_c_0), .B(SHAREDBUS_DAT_I[24]), .C(n29830), 
         .D(n34966), .Z(n36339)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i31167_4_lut.init = 16'hcaaa;
    LUT4 i31168_4_lut (.A(PIO_DATAI_adj_6643[0]), .B(LED_B_c_0), .C(n30231), 
         .D(n34926), .Z(n36340)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B+!(C (D))))) */ ;
    defparam i31168_4_lut.init = 16'h3aaa;
    CCU2C _add_1_add_4_16 (.A0(b[13]), .B0(p[12]), .C0(GND_net), .D0(VCC_net), 
          .A1(b[14]), .B1(p[13]), .C1(GND_net), .D1(VCC_net), .CIN(n27451), 
          .COUT(n27452), .S0(t[13]), .S1(t[14]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam _add_1_add_4_16.INIT0 = 16'h9995;
    defparam _add_1_add_4_16.INIT1 = 16'h9995;
    defparam _add_1_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_14 (.A0(b[11]), .B0(p[10]), .C0(GND_net), .D0(VCC_net), 
          .A1(b[12]), .B1(p[11]), .C1(GND_net), .D1(VCC_net), .CIN(n27450), 
          .COUT(n27451), .S0(t[11]), .S1(t[12]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam _add_1_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_12 (.A0(b[9]), .B0(p[8]), .C0(GND_net), .D0(VCC_net), 
          .A1(b[10]), .B1(p[9]), .C1(GND_net), .D1(VCC_net), .CIN(n27449), 
          .COUT(n27450), .S0(t[9]), .S1(t[10]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam _add_1_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_10 (.A0(b[7]), .B0(p[6]), .C0(GND_net), .D0(VCC_net), 
          .A1(b[8]), .B1(p[7]), .C1(GND_net), .D1(VCC_net), .CIN(n27448), 
          .COUT(n27449), .S0(t[7]), .S1(t[8]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam _add_1_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_8 (.A0(b[5]), .B0(p[4]), .C0(GND_net), .D0(VCC_net), 
          .A1(b[6]), .B1(p[5]), .C1(GND_net), .D1(VCC_net), .CIN(n27447), 
          .COUT(n27448), .S0(t[5]), .S1(t[6]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam _add_1_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_6 (.A0(b[3]), .B0(p[2]), .C0(GND_net), .D0(VCC_net), 
          .A1(b[4]), .B1(p[3]), .C1(GND_net), .D1(VCC_net), .CIN(n27446), 
          .COUT(n27447), .S0(t[3]), .S1(t[4]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam _add_1_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_4 (.A0(b[1]), .B0(p[0]), .C0(GND_net), .D0(VCC_net), 
          .A1(b[2]), .B1(p[1]), .C1(GND_net), .D1(VCC_net), .CIN(n27445), 
          .COUT(n27446), .S0(t[1]), .S1(t[2]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam _add_1_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_add_4_4.INJECT1_1 = "NO";
    PFUMX i33563 (.BLUT(n38964), .ALUT(n38963), .C0(LM32D_CYC_O), .Z(n38965));
    LUT4 i31163_3_lut_3_lut_4_lut (.A(write_idx_w[0]), .B(write_idx_w[1]), 
         .C(n6574), .D(n41325), .Z(n36335)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i31163_3_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i31158_3_lut_3_lut_4_lut (.A(write_idx_w[0]), .B(write_idx_w[1]), 
         .C(n6594), .D(n41325), .Z(n36330)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i31158_3_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i31153_3_lut_3_lut_4_lut (.A(write_idx_w[0]), .B(write_idx_w[1]), 
         .C(n6614), .D(n41325), .Z(n36325)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i31153_3_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i31149_3_lut_3_lut (.A(write_idx_w[0]), .B(write_idx_w[1]), .C(n6424), 
         .Z(n36321)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i31149_3_lut_3_lut.init = 16'hf1f1;
    LUT4 equal_2812_i2_1_lut_rep_1020 (.A(write_idx_w[4]), .Z(n41425)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam equal_2812_i2_1_lut_rep_1020.init = 16'h5555;
    LUT4 i3147_2_lut_4_lut_4_lut (.A(write_idx_w[4]), .B(counter[2]), .C(dcache_refill_request), 
         .D(n41430), .Z(n7610)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i3147_2_lut_4_lut_4_lut.init = 16'h0400;
    LUT4 i32068_3_lut (.A(n37237), .B(n37238), .C(write_idx_w[2]), .Z(n37240)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32068_3_lut.init = 16'hcaca;
    LUT4 i32067_3_lut (.A(n37235), .B(n37236), .C(write_idx_w[2]), .Z(n37239)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32067_3_lut.init = 16'hcaca;
    LUT4 i31161_3_lut_3_lut_4_lut (.A(write_idx_w[0]), .B(write_idx_w[1]), 
         .C(n6579), .D(n41325), .Z(n36333)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i31161_3_lut_3_lut_4_lut.init = 16'hf2f0;
    LUT4 i31157_3_lut_3_lut_4_lut (.A(write_idx_w[0]), .B(write_idx_w[1]), 
         .C(n6599), .D(n41325), .Z(n36329)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i31157_3_lut_3_lut_4_lut.init = 16'hf2f0;
    LUT4 i31148_3_lut_3_lut (.A(write_idx_w[0]), .B(write_idx_w[1]), .C(n6429), 
         .Z(n36320)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i31148_3_lut_3_lut.init = 16'hf2f2;
    LUT4 i31152_3_lut_3_lut_4_lut (.A(write_idx_w[0]), .B(write_idx_w[1]), 
         .C(n6619), .D(n41325), .Z(n36324)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i31152_3_lut_3_lut_4_lut.init = 16'hf2f0;
    LUT4 equal_2677_i6_2_lut_rep_1027 (.A(write_idx_w[2]), .B(write_idx_w[3]), 
         .Z(n41432)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam equal_2677_i6_2_lut_rep_1027.init = 16'heeee;
    LUT4 i31147_3_lut_3_lut (.A(write_idx_w[2]), .B(write_idx_w[3]), .C(n6439), 
         .Z(n36319)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i31147_3_lut_3_lut.init = 16'hf1f1;
    platform1_vhd inst_cpu (.\SHAREDBUS_ADR_I[7] (SHAREDBUS_ADR_I[7]), .n3(n3), 
            .\SHAREDBUS_ADR_I[10] (SHAREDBUS_ADR_I[10]), .n41347(n41347), 
            .n41303(n41303), .REF_CLK_c(REF_CLK_c), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .n41434(n41434), .inst1_FIFOof_wr(inst1_FIFOof_wr), .n41301(n41301), 
            .n41310(n41310), .inst3_Full(inst3_Full), .inst1_FIFOif_rd(inst1_FIFOif_rd), 
            .n35647(n35647), .inst3_Empty(inst3_Empty), .n41298(n41298), 
            .n41300(n41300), .n29(n29), .n41263(n41263), .\SHAREDBUS_ADR_I[29] (SHAREDBUS_ADR_I[29]), 
            .\SHAREDBUS_ADR_I[23] (SHAREDBUS_ADR_I[23]), .n45101(n45101), 
            .\counter[2] (counter[2]), .n12428(n12428), .n41346(n41346), 
            .n2(n2), .\selected[0] (selected[0]), .n32312(n32312), .\SHAREDBUS_ADR_I[5] (SHAREDBUS_ADR_I[5]), 
            .n34966(n34966), .n34926(n34926), .\SHAREDBUS_ADR_I[22] (SHAREDBUS_ADR_I[22]), 
            .n34242(n34242), .n41344(n41344), .n41299(n41299), .n30231(n30231), 
            .PIO_DATAI({PIO_DATAI_adj_6643}), .sclk_N_5010(sclk_N_5010), 
            .IO_SCK_c(IO_SCK_c), .rx_shift_data_31__N_4339(rx_shift_data_31__N_4339), 
            .n41328(n41328), .REF_CLK_c_enable_1453(REF_CLK_c_enable_1453), 
            .IO_MISO_c(IO_MISO_c), .IO_0_c_0(IO_0_c_0), .GND_net(GND_net), 
            .VCC_net(VCC_net), .IO_MOSI_c(IO_MOSI_c), .n41329(n41329), 
            .n41330(n41330), .n41331(n41331), .n41332(n41332), .n41333(n41333), 
            .n41334(n41334), .n41335(n41335), .\SHAREDBUS_DAT_I[8] (SHAREDBUS_DAT_I[8]), 
            .\SHAREDBUS_DAT_I[9] (SHAREDBUS_DAT_I[9]), .\SHAREDBUS_DAT_I[10] (SHAREDBUS_DAT_I[10]), 
            .\SHAREDBUS_DAT_I[11] (SHAREDBUS_DAT_I[11]), .\SHAREDBUS_DAT_I[12] (SHAREDBUS_DAT_I[12]), 
            .\SHAREDBUS_DAT_I[13] (SHAREDBUS_DAT_I[13]), .\SHAREDBUS_DAT_I[14] (SHAREDBUS_DAT_I[14]), 
            .\SHAREDBUS_DAT_I[15] (SHAREDBUS_DAT_I[15]), .n41336(n41336), 
            .n41337(n41337), .n41338(n41338), .n41339(n41339), .n41340(n41340), 
            .n41341(n41341), .n41342(n41342), .n41343(n41343), .\SHAREDBUS_DAT_I[24] (SHAREDBUS_DAT_I[24]), 
            .\SHAREDBUS_DAT_I[25] (SHAREDBUS_DAT_I[25]), .\SHAREDBUS_DAT_I[26] (SHAREDBUS_DAT_I[26]), 
            .\SHAREDBUS_DAT_I[27] (SHAREDBUS_DAT_I[27]), .\SHAREDBUS_DAT_I[28] (SHAREDBUS_DAT_I[28]), 
            .\SHAREDBUS_DAT_I[29] (SHAREDBUS_DAT_I[29]), .\SHAREDBUS_DAT_I[30] (SHAREDBUS_DAT_I[30]), 
            .\SHAREDBUS_DAT_I[31] (SHAREDBUS_DAT_I[31]), .n45179(n45179), 
            .n41380(n41380), .\inst_reg[15] (inst_reg[15]), .n10865(n10865), 
            .n41191(n41191), .\genblk1.read_address[10] (\genblk1.read_address [10]), 
            .\genblk1.write_address[10] (\genblk1.write_address [10]), .n3700(n3700), 
            .n5386(n5386), .n5085(n5085), .n3432(n3432), .\genblk1.state[2] (\genblk1.state [2]), 
            .\genblk1.pmi_address[3] (\genblk1.pmi_address [3]), .\genblk1.pmi_address[4] (\genblk1.pmi_address [4]), 
            .\genblk1.pmi_address[5] (\genblk1.pmi_address [5]), .\genblk1.pmi_address[6] (\genblk1.pmi_address [6]), 
            .\genblk1.pmi_address[7] (\genblk1.pmi_address [7]), .\genblk1.pmi_address[8] (\genblk1.pmi_address [8]), 
            .\genblk1.pmi_address[9] (\genblk1.pmi_address [9]), .\genblk1.pmi_address[10] (\genblk1.pmi_address [10]), 
            .\genblk1.pmi_address[11] (\genblk1.pmi_address [11]), .\genblk1.pmi_address[12] (\genblk1.pmi_address [12]), 
            .\genblk1.pmi_address[13] (\genblk1.pmi_address [13]), .\genblk1.pmi_address[14] (\genblk1.pmi_address [14]), 
            .n41321(n41321), .n20000(n20000), .n6038(n6038), .n11843(n11843), 
            .n3485(n3485), .n6034(n6034), .n41292(n41292), .n19822(n19822), 
            .n41390(n41390), .n3486(n3486), .n82_adj_343({n34_adj_6597, 
            n37_adj_6598, n40, n43, n46, n49, n52, n55, n58, 
            n61, n64_adj_6599, n67_adj_6600, n70_adj_6601, n73_adj_6602, 
            n76_adj_6603}), .n45076(n45076), .n8(n8), .LM32D_CYC_O(LM32D_CYC_O), 
            .locked_N_493(locked_N_493), .\LM32D_CTI_O[0] (LM32D_CTI_O[0]), 
            .\LM32I_ADR_O[12] (LM32I_ADR_O[12]), .n29830(n29830), .\next_cycle_type[2] (next_cycle_type_adj_6725[2]), 
            .write_idx_w({write_idx_w}), .n41352(n41352), .n41351(n41351), 
            .w_result({w_result}), .n41350(n41350), .dcache_refill_request(dcache_refill_request), 
            .\operand_1_x[1] (operand_1_x[1]), .dc_re(dc_re), .n41430(n41430), 
            .n41432(n41432), .REF_CLK_c_enable_176(REF_CLK_c_enable_176), 
            .n7611(n7611), .n41405(n41405), .REF_CLK_c_enable_164(REF_CLK_c_enable_164), 
            .n41356(n41356), .n41355(n41355), .n41353(n41353), .n41358(n41358), 
            .n41359(n41359), .\operand_m[10] (operand_m[10]), .\operand_m[9] (operand_m[9]), 
            .\operand_m[5] (operand_m[5]), .dcache_select_x(dcache_select_x), 
            .n41354(n41354), .bie(bie), .n31279(n31279), .\adder_result_x[16] (adder_result_x[16]), 
            .\adder_result_x[17] (adder_result_x[17]), .\adder_result_x[18] (adder_result_x[18]), 
            .\adder_result_x[19] (adder_result_x[19]), .\adder_result_x[20] (adder_result_x[20]), 
            .\adder_result_x[21] (adder_result_x[21]), .\adder_result_x[22] (adder_result_x[22]), 
            .\adder_result_x[23] (adder_result_x[23]), .\adder_result_x[24] (adder_result_x[24]), 
            .\adder_result_x[25] (adder_result_x[25]), .\adder_result_x[26] (adder_result_x[26]), 
            .\adder_result_x[27] (adder_result_x[27]), .\adder_result_x[28] (adder_result_x[28]), 
            .\adder_result_x[29] (adder_result_x[29]), .\adder_result_x[30] (adder_result_x[30]), 
            .\adder_result_x[31] (adder_result_x[31]), .n6518(n6518), .n6648(n6648), 
            .branch_target_d({branch_target_d}), .direction_m(direction_m), 
            .n45103(n45103), .n45099(n45099), .n41394(n41394), .n41401(n41401), 
            .bie_N_3274(bie_N_3274), .pc_f({pc_f}), .n41325(n41325), .n17816(n17816), 
            .n41379(n41379), .\shifter_result_m[21] (shifter_result_m[21]), 
            .n41357(n41357), .\left_shift_result[21] (left_shift_result[21]), 
            .\left_shift_result[10] (left_shift_result[10]), .b({b}), .\p[0] (p[0]), 
            .\p[1] (p[1]), .\p[2] (p[2]), .\p[3] (p[3]), .\p[4] (p[4]), 
            .\p[5] (p[5]), .\p[6] (p[6]), .\p[7] (p[7]), .\p[8] (p[8]), 
            .\p[9] (p[9]), .\p[10] (p[10]), .\p[11] (p[11]), .\p[12] (p[12]), 
            .\p[13] (p[13]), .\p[14] (p[14]), .\p[15] (p[15]), .\p[16] (p[16]), 
            .\p[17] (p[17]), .\p[18] (p[18]), .\p[19] (p[19]), .\p[20] (p[20]), 
            .\p[21] (p[21]), .\p[22] (p[22]), .\p[23] (p[23]), .\p[24] (p[24]), 
            .\p[25] (p[25]), .\p[26] (p[26]), .\p[27] (p[27]), .\p[28] (p[28]), 
            .\p[29] (p[29]), .\p[30] (p[30]), .\a[31] (a[31]), .t({t}), 
            .n38965(n38965), .\d_adr_o_31__N_2278[5] (d_adr_o_31__N_2278[5]), 
            .\d_adr_o_31__N_2278[9] (d_adr_o_31__N_2278[9]), .\d_adr_o_31__N_2278[10] (d_adr_o_31__N_2278[10]), 
            .\LM32D_ADR_O[17] (LM32D_ADR_O[17]), .\LM32D_ADR_O[19] (LM32D_ADR_O[19]), 
            .\state[0] (state_adj_6798[0]), .\state[2] (state_adj_6798[2]), 
            .flush_set({flush_set_adj_6801}), .flush_set_8__N_2513({flush_set_8__N_2513}), 
            .\dcache_refill_address[5] (dcache_refill_address[5]), .\dcache_refill_address[9] (dcache_refill_address[9]), 
            .\dcache_refill_address[10] (dcache_refill_address[10]), .\tmem_write_address[1] (tmem_write_address_adj_6794[1]), 
            .\tmem_write_address[5] (tmem_write_address_adj_6794[5]), .\tmem_write_address[6] (tmem_write_address_adj_6794[6]), 
            .\dmem_write_address[3] (dmem_write_address_adj_6796[3]), .\dmem_write_address[7] (dmem_write_address_adj_6796[7]), 
            .\dmem_write_address[8] (dmem_write_address_adj_6796[8]), .n36337(n36337), 
            .n6781(n6781), .n6764(n6764), .n6749(n6749), .pc_d({pc_d}), 
            .n6760(n6760), .n45105(n45105), .n6589(n6589), .n6584(n6584), 
            .n37179(n37179), .n6439(n6439), .n6434(n6434), .n37177(n37177), 
            .n6599(n6599), .n6594(n6594), .n37180(n37180), .n6629(n6629), 
            .n6624(n6624), .n37183(n37183), .n6579(n6579), .n6574(n6574), 
            .n37178(n37178), .n6429(n6429), .n6424(n6424), .n37176(n37176), 
            .n6609(n6609), .n6604(n6604), .n37181(n37181), .n6619(n6619), 
            .n6614(n6614), .n37182(n37182), .n37185(n37185), .n37184(n37184), 
            .n37188(n37188), .n37187(n37187), .n37186(n37186), .n37189(n37189), 
            .n7603(n7603), .n7571(n7571), .n7607(n7607), .n7575(n7575), 
            .n7606(n7606), .n7574(n7574), .n7604(n7604), .n7572(n7572), 
            .n7605(n7605), .n7573(n7573), .n7608(n7608), .n7576(n7576), 
            .n7602(n7602), .n7570(n7570), .n7601(n7601), .n7569(n7569), 
            .n7600(n7600), .n7568(n7568), .n7599(n7599), .n7567(n7567), 
            .n7598(n7598), .n7566(n7566), .n7597(n7597), .n7565(n7565), 
            .n7596(n7596), .n7564(n7564), .n7595(n7595), .n7563(n7563), 
            .n7594(n7594), .n7562(n7562), .n7593(n7593), .n7561(n7561), 
            .n7592(n7592), .n7560(n7560), .n7584(n7584), .n7552(n7552), 
            .n7583(n7583), .n7551(n7551), .n7582(n7582), .n7550(n7550), 
            .n7581(n7581), .n7549(n7549), .n7580(n7580), .n7548(n7548), 
            .n7579(n7579), .n7547(n7547), .n7578(n7578), .n7546(n7546), 
            .n7577(n7577), .n7545(n7545), .n6750(n6750), .n7591(n7591), 
            .n7559(n7559), .n7590(n7590), .n7558(n7558), .n7589(n7589), 
            .n7557(n7557), .n7588(n7588), .n7556(n7556), .n7587(n7587), 
            .n7555(n7555), .n7586(n7586), .n7554(n7554), .n7585(n7585), 
            .n7553(n7553), .n37501(n37501), .n37500(n37500), .n37502(n37502), 
            .n37499(n37499), .n37498(n37498), .n37497(n37497), .n37496(n37496), 
            .n6751(n6751), .n6752(n6752), .n6753(n6753), .n6754(n6754), 
            .n6755(n6755), .n6756(n6756), .n6757(n6757), .n6758(n6758), 
            .n6759(n6759), .n6761(n6761), .n6762(n6762), .n6763(n6763), 
            .n37495(n37495), .n7672(n7672), .n7640(n7640), .n7673(n7673), 
            .n7641(n7641), .n34_adj_327(n34), .n7674(n7674), .n7642(n7642), 
            .n7675(n7675), .n7643(n7643), .n7676(n7676), .n7644(n7644), 
            .n7671(n7671), .n7639(n7639), .n7670(n7670), .n7638(n7638), 
            .n7669(n7669), .n7637(n7637), .n7668(n7668), .n7636(n7636), 
            .n7667(n7667), .n7635(n7635), .n7666(n7666), .n7634(n7634), 
            .n7665(n7665), .n7633(n7633), .n7664(n7664), .n7632(n7632), 
            .n7663(n7663), .n7631(n7631), .n7662(n7662), .n7630(n7630), 
            .n7661(n7661), .n7629(n7629), .n7660(n7660), .n7628(n7628), 
            .n36(n36), .n7652(n7652), .n7620(n7620), .n7651(n7651), 
            .n7619(n7619), .n7650(n7650), .n7618(n7618), .n7649(n7649), 
            .n7617(n7617), .n37_adj_328(n37), .n7648(n7648), .n7616(n7616), 
            .n7647(n7647), .n7615(n7615), .n7646(n7646), .n7614(n7614), 
            .n7645(n7645), .n7613(n7613), .n7659(n7659), .n7627(n7627), 
            .n7658(n7658), .n7626(n7626), .n7657(n7657), .n7625(n7625), 
            .n7656(n7656), .n7624(n7624), .n7655(n7655), .n7623(n7623), 
            .n7654(n7654), .n7622(n7622), .n7653(n7653), .n7621(n7621), 
            .n37504(n37504), .n37503(n37503), .n37507(n37507), .n37506(n37506), 
            .n37505(n37505), .n37508(n37508), .n45106(n45106), .\LM32I_ADR_O[17] (LM32I_ADR_O[17]), 
            .\LM32I_ADR_O[19] (LM32I_ADR_O[19]), .flush_set_adj_344({flush_set}), 
            .flush_set_8__N_1953({flush_set_8__N_1953}), .n157({n64, n67, 
            n70, n73, n76, n79, n82, n85, n88, n91, n94, n97, 
            n100, n103, n106, n109, n112, n115, n118, n121, 
            n124, n127, n130, n133, n136, n139, n142, n145, 
            n148, n151}), .n36336(n36336), .n10589(n10589), .n10585(n10585), 
            .n10591(n10591), .n10593(n10593), .n10587(n10587), .n10595(n10595), 
            .n10452(n10452), .LED_R_c_0(LED_R_c_0), .n36338(n36338), .LED_G_c_0(LED_G_c_0), 
            .LED_B_c_0(LED_B_c_0), .n36339(n36339), .n36340(n36340), .n35006(n35006), 
            .inst1_FIFOfifo_rst(inst1_FIFOfifo_rst), .inst3_Q({inst3_Q}));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(86[12:37])
    LUT4 i12499_3_lut (.A(left_shift_result[21]), .B(left_shift_result[10]), 
         .C(direction_m), .Z(n17816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(92[5:16])
    defparam i12499_3_lut.init = 16'hcaca;
    LUT4 i12519_3_lut (.A(left_shift_result[10]), .B(left_shift_result[21]), 
         .C(direction_m), .Z(shifter_result_m[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(92[5:16])
    defparam i12519_3_lut.init = 16'hcaca;
    fifo_dc_32x32 inst3 (.inst3_Full(inst3_Full), .REF_CLK_c(REF_CLK_c), 
            .inst1_FIFOfifo_rst(inst1_FIFOfifo_rst), .inst3_Empty(inst3_Empty), 
            .GND_net(GND_net), .VCC_net(VCC_net), .inst1_FIFOof_wr(inst1_FIFOof_wr), 
            .inst1_FIFOif_rd(inst1_FIFOif_rd), .\SHAREDBUS_DAT_I[31] (SHAREDBUS_DAT_I[31]), 
            .\SHAREDBUS_DAT_I[30] (SHAREDBUS_DAT_I[30]), .\SHAREDBUS_DAT_I[29] (SHAREDBUS_DAT_I[29]), 
            .\SHAREDBUS_DAT_I[28] (SHAREDBUS_DAT_I[28]), .\SHAREDBUS_DAT_I[27] (SHAREDBUS_DAT_I[27]), 
            .\SHAREDBUS_DAT_I[26] (SHAREDBUS_DAT_I[26]), .\SHAREDBUS_DAT_I[25] (SHAREDBUS_DAT_I[25]), 
            .\SHAREDBUS_DAT_I[24] (SHAREDBUS_DAT_I[24]), .n41343(n41343), 
            .n41342(n41342), .n41341(n41341), .n41340(n41340), .n41339(n41339), 
            .n41338(n41338), .n41337(n41337), .n41336(n41336), .\SHAREDBUS_DAT_I[15] (SHAREDBUS_DAT_I[15]), 
            .\SHAREDBUS_DAT_I[14] (SHAREDBUS_DAT_I[14]), .\SHAREDBUS_DAT_I[13] (SHAREDBUS_DAT_I[13]), 
            .\SHAREDBUS_DAT_I[12] (SHAREDBUS_DAT_I[12]), .\SHAREDBUS_DAT_I[11] (SHAREDBUS_DAT_I[11]), 
            .\SHAREDBUS_DAT_I[10] (SHAREDBUS_DAT_I[10]), .\SHAREDBUS_DAT_I[9] (SHAREDBUS_DAT_I[9]), 
            .\SHAREDBUS_DAT_I[8] (SHAREDBUS_DAT_I[8]), .n41335(n41335), 
            .n41334(n41334), .n41333(n41333), .n41332(n41332), .n41331(n41331), 
            .n41330(n41330), .n41329(n41329), .n41328(n41328), .inst3_Q({inst3_Q})) /* synthesis NGD_DRC_MASK=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    LUT4 m0_lut (.Z(n45086)) /* synthesis lut_function=0, syn_instantiated=1 */ ;
    defparam m0_lut.init = 16'h0000;
    VLO i1 (.Z(GND_net));
    PFUMX i32018 (.BLUT(n37188), .ALUT(n37189), .C0(n41353), .Z(n37190));
    LUT4 i2824_4_lut (.A(n6642), .B(n37509), .C(n6645), .D(n41357), 
         .Z(n6648)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i2824_4_lut.init = 16'hc088;
    
endmodule
//
// Verilog Description of module fpgacfg
//

module fpgacfg (sclk_N_5010, n41434, VCC_net, \from_fpgacfg.wfm_ch_en , 
            REF_CLK_c, \from_fpgacfg.CLK_ENA , IO_MOSI_c, \from_fpgacfg.FX3_LED_CTRL , 
            \from_fpgacfg.FPGA_LED1_CTRL , \from_fpgacfg.GPIO , \from_fpgacfg.txant_post , 
            \from_fpgacfg.txant_pre , \from_fpgacfg.sync_size , \inst2_from_fpgacfg.wfm_smpl_width[0] , 
            \inst2_from_fpgacfg.rx_en , \inst2_from_fpgacfg.smpl_nr_clr , 
            \from_fpgacfg.smpl_width , \from_fpgacfg.ch_en , \from_fpgacfg.clk_ind , 
            \from_fpgacfg.drct_clk_en , \from_fpgacfg.phase_reg_sel , IO_0_c_0, 
            \from_fpgacfg.SPI_SS , \inst2_from_fpgacfg.load_phase_reg , 
            \inst2_from_fpgacfg.synch_mode , \inst2_from_fpgacfg.tx_cnt_en , 
            \from_fpgacfg.sync_pulse_period , \inst2_from_fpgacfg.wfm_load , 
            \inst2_from_fpgacfg.wfm_play , REF_CLK_c_enable_1424, \inst2_from_fpgacfg.LMS1_RXEN , 
            \inst2_from_fpgacfg.LMS1_TXEN , \inst2_from_fpgacfg.LMS1_TXNRX2 , 
            \inst2_from_fpgacfg.LMS1_TXNRX1 , \inst2_from_fpgacfg.LMS1_CORE_LDO_EN , 
            \inst2_from_fpgacfg.LMS1_RESET , \from_fpgacfg.FPGA_LED2_CTRL , 
            \inst2_from_fpgacfg.LMS1_SS , \inst2_from_fpgacfg.tx_en , \inst2_from_fpgacfg.rx_ptrn_en , 
            \inst2_from_fpgacfg.tx_ptrn_en , \inst2_from_fpgacfg.txpct_loss_clr , 
            \inst2_from_fpgacfg.mode , \inst2_from_fpgacfg.ddr_en , \inst2_from_fpgacfg.trxiq_pulse , 
            \inst2_from_fpgacfg.mimo_int_en , \inst2_from_fpgacfg.synch_dis , 
            \from_fpgacfg.cnt_ind , n41191, \inst_reg[15] , REF_CLK_c_enable_1453, 
            n45086, n10865, n2023, rx_shift_data_31__N_4339, IO_MISO_c, 
            n45179, n35448, USER_BUTTON_c);
    input sclk_N_5010;
    output n41434;
    input VCC_net;
    output [15:0]\from_fpgacfg.wfm_ch_en ;
    input REF_CLK_c;
    output [3:0]\from_fpgacfg.CLK_ENA ;
    input IO_MOSI_c;
    output [2:0]\from_fpgacfg.FX3_LED_CTRL ;
    output [2:0]\from_fpgacfg.FPGA_LED1_CTRL ;
    output [15:0]\from_fpgacfg.GPIO ;
    output [15:0]\from_fpgacfg.txant_post ;
    output [15:0]\from_fpgacfg.txant_pre ;
    output [15:0]\from_fpgacfg.sync_size ;
    output \inst2_from_fpgacfg.wfm_smpl_width[0] ;
    output \inst2_from_fpgacfg.rx_en ;
    output \inst2_from_fpgacfg.smpl_nr_clr ;
    output [1:0]\from_fpgacfg.smpl_width ;
    output [15:0]\from_fpgacfg.ch_en ;
    output [4:0]\from_fpgacfg.clk_ind ;
    output [15:0]\from_fpgacfg.drct_clk_en ;
    output [15:0]\from_fpgacfg.phase_reg_sel ;
    input IO_0_c_0;
    output [15:0]\from_fpgacfg.SPI_SS ;
    output \inst2_from_fpgacfg.load_phase_reg ;
    output \inst2_from_fpgacfg.synch_mode ;
    output \inst2_from_fpgacfg.tx_cnt_en ;
    output [31:0]\from_fpgacfg.sync_pulse_period ;
    output \inst2_from_fpgacfg.wfm_load ;
    output \inst2_from_fpgacfg.wfm_play ;
    input REF_CLK_c_enable_1424;
    output \inst2_from_fpgacfg.LMS1_RXEN ;
    output \inst2_from_fpgacfg.LMS1_TXEN ;
    output \inst2_from_fpgacfg.LMS1_TXNRX2 ;
    output \inst2_from_fpgacfg.LMS1_TXNRX1 ;
    output \inst2_from_fpgacfg.LMS1_CORE_LDO_EN ;
    output \inst2_from_fpgacfg.LMS1_RESET ;
    output [2:0]\from_fpgacfg.FPGA_LED2_CTRL ;
    output \inst2_from_fpgacfg.LMS1_SS ;
    output \inst2_from_fpgacfg.tx_en ;
    output \inst2_from_fpgacfg.rx_ptrn_en ;
    output \inst2_from_fpgacfg.tx_ptrn_en ;
    output \inst2_from_fpgacfg.txpct_loss_clr ;
    output \inst2_from_fpgacfg.mode ;
    output \inst2_from_fpgacfg.ddr_en ;
    output \inst2_from_fpgacfg.trxiq_pulse ;
    output \inst2_from_fpgacfg.mimo_int_en ;
    output \inst2_from_fpgacfg.synch_dis ;
    output [4:0]\from_fpgacfg.cnt_ind ;
    input n41191;
    output \inst_reg[15] ;
    input REF_CLK_c_enable_1453;
    input n45086;
    output n10865;
    output n2023;
    input rx_shift_data_31__N_4339;
    output IO_MISO_c;
    input n45179;
    output n35448;
    input USER_BUTTON_c;
    
    wire sclk_N_5010 /* synthesis is_inv_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(57[11:19])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire [15:0]dout_reg;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(57[11:19])
    
    wire sclk_N_5010_enable_16;
    wire [15:0]dout_reg_15__N_4993;
    wire [3:0]hw_ver_int;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(66[11:21])
    wire [15:0]\mem[3] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    wire [15:0]\mem[2] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    wire [15:0]inst_reg;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(51[11:19])
    
    wire n37363, REF_CLK_c_enable_205;
    wire [15:0]din_reg;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(54[11:18])
    
    wire REF_CLK_c_enable_387, REF_CLK_c_enable_384;
    wire [15:0]\mem[27] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    
    wire REF_CLK_c_enable_382;
    wire [15:0]\mem[9] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    wire [15:0]\mem[8] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    
    wire n37315;
    wire [15:0]\mem[11] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    wire [15:0]\mem[10] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    
    wire n37314;
    wire [15:0]\mem[13] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    
    wire n37313, REF_CLK_c_enable_367;
    wire [15:0]\mem[25] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    
    wire REF_CLK_c_enable_352;
    wire [15:0]\mem[24] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    
    wire REF_CLK_c_enable_337, REF_CLK_c_enable_322;
    wire [15:0]\mem[22] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    
    wire REF_CLK_c_enable_304;
    wire [15:0]\mem[21] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    
    wire REF_CLK_c_enable_289;
    wire [15:0]\mem[20] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    
    wire REF_CLK_c_enable_273;
    wire [15:0]\mem[19] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    
    wire REF_CLK_c_enable_258;
    wire [15:0]\mem[18] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    
    wire REF_CLK_c_enable_242, REF_CLK_c_enable_226, REF_CLK_c_enable_211, 
        REF_CLK_c_enable_174;
    wire [15:0]\mem[14] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    
    wire REF_CLK_c_enable_119, REF_CLK_c_enable_101, REF_CLK_c_enable_511, 
        REF_CLK_c_enable_526, REF_CLK_c_enable_541, REF_CLK_c_enable_556, 
        REF_CLK_c_enable_571, REF_CLK_c_enable_586, REF_CLK_c_enable_601, 
        REF_CLK_c_enable_616, REF_CLK_c_enable_631, REF_CLK_c_enable_646;
    wire [15:0]\mem[1] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    
    wire REF_CLK_c_enable_661;
    wire [15:0]\mem[0] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    
    wire REF_CLK_c_enable_676, n37312, n26, n27, n37480, n37308, 
        n37362, n37361, n37307, n37357, n37356, n37306, n37305, 
        n37301, n37300, n37299, n31786;
    wire [15:0]\mem[6] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    
    wire n37298, n37294, n37293, n37292, n37291, n37287, n37286, 
        REF_CLK_c_enable_202, n37285, n37284, REF_CLK_c_enable_1608, 
        n37355, n37354, n37350, n37349, n37280, n37279, n37278, 
        n37348, n37347, n37277, n37343, n37342, n37341, n37273, 
        n37340, n37272, n37271, n37270;
    wire [63:0]n1800;
    
    wire n11745, n41219, n37266, n37265, n37264, n37263, n37259, 
        n37258, n37257, n37256, n37252, n37336, n37251, n37250, 
        n37335, n37249, n37245, n37334, n37333, n37244, n37329, 
        n37328, n37243, n37242, n37327, n37326, n37322, n37321, 
        n37320, n37319, n41456, n41457, n41458, n36314;
    wire [15:0]\mem[26] ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(60[11:14])
    
    wire n36313, n41453, n41454, n41455, n37318, n37325, n35957, 
        n37339, n37346, n36011, n37360, n37367, n36026, n37255, 
        n37262, n36275, n37381, n37388, n36287, n37402, n37409, 
        n36290, n37193, n37194, n37196, n37465, n37472, n36050, 
        n37200, n37201, n37203, n37423, n37430, n36296, n37444, 
        n37451, n36299, n37207, n37208, n37210, n37276, n37283, 
        n36302, n37297, n37304, n36311, n37483, n37484, n37486, 
        n37490, n37491, n37493, n35985, n35988, n37192, n35991, 
        n35994, n35997, n36000, n36006, n36009, n37199, n36015, 
        n36018, n36021, n36024, n36033, n36036, n37206, REF_CLK_c_enable_1621, 
        n36039, n36042, n36045, n36048, n37246, n37247, n37248, 
        n37253, n37254, n37260, n37261, n37267, n37268, n37269, 
        n37274, n37275, n37281, n37282, n37288, n37289, n37290, 
        n37295, n37296, n37302, n37303, n37309, n37310, n37311, 
        n37316, n37317, n37323, n37324, n37330, n37331, n37332, 
        n37337, n37338, n37344, n37345, n37351, n37352, n37353, 
        n36308, n37358, n37359, n37365, n37366, n37372, n37373, 
        n37374, n37379, n37380, n37386, n37387, n37393, n37394, 
        n37395, n37400, n37401, n37407, n37408, n37414, n37415, 
        n37416, n37421, n37422, n36307, n37428, n37429, n37435, 
        n37436, n37437, n37442, n37443, n37449, n37450, n37456, 
        n37457, n37458, n36305, n37463, n37464, n37470, n37471, 
        n37473, n37474, n37481, n36304, n36293, n36292, n37475, 
        n37476, n37482, n37477, n37478, n37479, n36168, n36165, 
        n37489, n36162, n36159, n36156, n36153, n36047, n36046, 
        n36044, n37492;
    wire [15:0]dout_reg_15__N_5274;
    
    wire n36043, n36041, n36040, n36038, n36037, n36035, n36034, 
        n36032, n36031, n37488, n41431, n36174, n36023, n36022, 
        n37195, n37191, n20513, n35982, n37202, n37485, n36020, 
        n36019, n36017, n37209, n36016, n11789, n41446, n30140, 
        n31780, n30139, n11264, n24, n41384, n35959, n35960, n35961, 
        n41447, n35962, n35963, n35964, n23, n41174, n36294, n36274, 
        n36306, n36301, n36309, n36310, n36315, n35956, n36010, 
        n36025, n35967, n36286, n35965, n35966, n35970, n36289, 
        n35973, n36295, n35976, n36298, n35979, n36049, n35968, 
        n35969, n35971, n35972, n35974, n35975, n35977, n35978, 
        n20, n19, n17, n35980, n35981, n35983, n35984, n36014, 
        n35986, n35987, n35989, n35990, n35992, n35993, n35995, 
        n35996, n35998, n35999, n36013, n36008, n16, n12, n36004, 
        n36005, n36007, n11, n9, n8, n5, n4, n36173, n36172, 
        n36167, n36166, n36164, n36163, n37469, n37468, n37467, 
        n37466, n36161, n36160, n36158, n36157, n36155, n36154, 
        n36152, n36151, n37462, n37461, n37460, n37459, n37455, 
        n37454, n37453, n37452, n37448, n37447, n37446, n37445, 
        n37441, n37440, n37439, n37438, n37434, n37433, n37432, 
        n37431, n37427, n37426, n41182, n41443, n37425, n37424, 
        n37420, n37419, n37418, n37417, n37413, n37412, n37411, 
        n37410, n37406, n37405, n37404, n37403, n37399, n37398, 
        n37397, n37396, n37392, n37391, n37390, n37389, n37364, 
        n37368, n37369, n37370, n37371, n37375, n37376, n37377, 
        n37378, n37382, n37383, n37384, n37385, n37957, n37958, 
        n36453;
    
    FD1P3DX dout_reg_i0 (.D(dout_reg_15__N_4993[0]), .SP(sclk_N_5010_enable_16), 
            .CK(sclk_N_5010), .CD(n41434), .Q(dout_reg[0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(151[7] 170[14])
    defparam dout_reg_i0.GSR = "ENABLED";
    FD1S3DX hw_ver_int_i1 (.D(VCC_net), .CK(sclk_N_5010), .CD(n41434), 
            .Q(hw_ver_int[2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(187[7] 202[14])
    defparam hw_ver_int_i1.GSR = "ENABLED";
    LUT4 i32191_3_lut (.A(\mem[3] [10]), .B(\mem[2] [10]), .C(inst_reg[0]), 
         .Z(n37363)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32191_3_lut.init = 16'hcaca;
    FD1P3DX mem_12__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_205), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.wfm_ch_en [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_12__i0_i10.GSR = "ENABLED";
    FD1P3BX mem_29__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_387), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.CLK_ENA [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_29__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_28__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_384), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.FX3_LED_CTRL [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_28__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_27__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_382), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[27] [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_27__i0_i0.GSR = "ENABLED";
    LUT4 i32143_3_lut (.A(\mem[9] [12]), .B(\mem[8] [12]), .C(inst_reg[0]), 
         .Z(n37315)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32143_3_lut.init = 16'hcaca;
    LUT4 i32142_3_lut (.A(\mem[11] [12]), .B(\mem[10] [12]), .C(inst_reg[0]), 
         .Z(n37314)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32142_3_lut.init = 16'hcaca;
    LUT4 i32141_3_lut (.A(\mem[13] [12]), .B(\from_fpgacfg.wfm_ch_en [12]), 
         .C(inst_reg[0]), .Z(n37313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32141_3_lut.init = 16'hcaca;
    FD1P3DX mem_26___i1 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_367), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.FPGA_LED1_CTRL [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_26___i1.GSR = "ENABLED";
    FD1P3DX mem_25__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_352), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[25] [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_25__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_24__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_337), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[24] [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_24__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_23__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_322), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.GPIO [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_23__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_22__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_304), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[22] [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_22__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_21__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_289), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[21] [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_21__i0_i0.GSR = "ENABLED";
    FD1P3BX mem_20__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_273), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[20] [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_20__i0_i0.GSR = "ENABLED";
    FD1P3BX mem_19__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_258), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[19] [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_19__i0_i0.GSR = "ENABLED";
    FD1P3BX mem_18__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_242), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[18] [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_18__i0_i0.GSR = "ENABLED";
    FD1P3BX mem_17__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_226), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.txant_post [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_17__i0_i0.GSR = "ENABLED";
    FD1P3BX mem_16__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_211), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.txant_pre [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_16__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_15__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_174), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_size [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_15__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_14__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_119), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[14] [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_14__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_13___i1 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_101), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\inst2_from_fpgacfg.wfm_smpl_width[0] )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_13___i1.GSR = "ENABLED";
    FD1P3BX mem_12__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_205), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.wfm_ch_en [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_12__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_11__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_511), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[11] [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_11__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_10___i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_526), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\inst2_from_fpgacfg.rx_en )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_10___i0.GSR = "ENABLED";
    FD1P3BX mem_9___i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_541), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\inst2_from_fpgacfg.smpl_nr_clr )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_9___i0.GSR = "ENABLED";
    FD1P3DX mem_8___i1 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_556), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.smpl_width [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_8___i1.GSR = "ENABLED";
    FD1P3BX mem_7__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_571), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.ch_en [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_7__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_6___i1 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_586), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.clk_ind [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_6___i1.GSR = "ENABLED";
    FD1P3DX mem_5__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_601), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.drct_clk_en [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_5__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_4__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_616), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.phase_reg_sel [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_4__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_3__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_631), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[3] [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_3__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_2__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_646), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[2] [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_2__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_1__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_661), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[1] [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_1__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_0__i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_676), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[0] [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_0__i0_i0.GSR = "ENABLED";
    FD1P3DX mem_12__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_205), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.wfm_ch_en [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_12__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_12__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_205), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.wfm_ch_en [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_12__i0_i8.GSR = "ENABLED";
    LUT4 i32140_3_lut (.A(\from_fpgacfg.sync_size [12]), .B(\mem[14] [12]), 
         .C(inst_reg[0]), .Z(n37312)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32140_3_lut.init = 16'hcaca;
    PFUMX i32308 (.BLUT(n26), .ALUT(n27), .C0(inst_reg[1]), .Z(n37480));
    LUT4 mem_18__15__I_0_207_i9_2_lut (.A(\mem[18] [8]), .B(IO_0_c_0), .Z(\from_fpgacfg.SPI_SS [8])) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(301[35:58])
    defparam mem_18__15__I_0_207_i9_2_lut.init = 16'hbbbb;
    FD1P3DX mem_12__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_205), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.wfm_ch_en [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_12__i0_i7.GSR = "ENABLED";
    LUT4 i32136_3_lut (.A(\from_fpgacfg.txant_post [12]), .B(\from_fpgacfg.txant_pre [12]), 
         .C(inst_reg[0]), .Z(n37308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32136_3_lut.init = 16'hcaca;
    FD1P3DX mem_12__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_205), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.wfm_ch_en [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_12__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_12__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_205), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.wfm_ch_en [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_12__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_12__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_205), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.wfm_ch_en [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_12__i0_i4.GSR = "ENABLED";
    LUT4 i32190_3_lut (.A(\from_fpgacfg.drct_clk_en [10]), .B(\from_fpgacfg.phase_reg_sel [10]), 
         .C(inst_reg[0]), .Z(n37362)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32190_3_lut.init = 16'hcaca;
    LUT4 i32189_3_lut (.A(\from_fpgacfg.ch_en [10]), .B(\inst2_from_fpgacfg.load_phase_reg ), 
         .C(inst_reg[0]), .Z(n37361)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32189_3_lut.init = 16'hcaca;
    LUT4 i32135_3_lut (.A(\mem[19] [12]), .B(\mem[18] [12]), .C(inst_reg[0]), 
         .Z(n37307)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32135_3_lut.init = 16'hcaca;
    LUT4 i32185_3_lut (.A(\mem[9] [10]), .B(\inst2_from_fpgacfg.synch_mode ), 
         .C(inst_reg[0]), .Z(n37357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32185_3_lut.init = 16'hcaca;
    LUT4 i32184_3_lut (.A(\mem[11] [10]), .B(\inst2_from_fpgacfg.tx_cnt_en ), 
         .C(inst_reg[0]), .Z(n37356)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32184_3_lut.init = 16'hcaca;
    LUT4 i32134_3_lut (.A(\mem[21] [12]), .B(\mem[20] [12]), .C(inst_reg[0]), 
         .Z(n37306)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32134_3_lut.init = 16'hcaca;
    LUT4 i32133_3_lut (.A(\from_fpgacfg.GPIO [12]), .B(\mem[22] [12]), .C(inst_reg[0]), 
         .Z(n37305)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32133_3_lut.init = 16'hcaca;
    LUT4 i32129_3_lut (.A(\mem[1] [13]), .B(\mem[0] [13]), .C(inst_reg[0]), 
         .Z(n37301)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32129_3_lut.init = 16'hcaca;
    LUT4 i32128_3_lut (.A(\mem[3] [13]), .B(\mem[2] [13]), .C(inst_reg[0]), 
         .Z(n37300)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32128_3_lut.init = 16'hcaca;
    LUT4 i32127_3_lut (.A(\from_fpgacfg.drct_clk_en [13]), .B(\from_fpgacfg.phase_reg_sel [13]), 
         .C(inst_reg[0]), .Z(n37299)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32127_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut (.A(inst_reg[2]), .B(inst_reg[3]), .C(inst_reg[4]), 
         .Z(n31786)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(253[20:62])
    defparam i1_3_lut.init = 16'hfbfb;
    LUT4 mem_18__15__I_0_207_i8_2_lut (.A(\mem[18] [7]), .B(IO_0_c_0), .Z(\from_fpgacfg.SPI_SS [7])) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(301[35:58])
    defparam mem_18__15__I_0_207_i8_2_lut.init = 16'hbbbb;
    LUT4 i32126_3_lut (.A(\from_fpgacfg.ch_en [13]), .B(\mem[6] [13]), .C(inst_reg[0]), 
         .Z(n37298)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32126_3_lut.init = 16'hcaca;
    LUT4 i32122_3_lut (.A(\mem[9] [13]), .B(\mem[8] [13]), .C(inst_reg[0]), 
         .Z(n37294)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32122_3_lut.init = 16'hcaca;
    LUT4 i32121_3_lut (.A(\mem[11] [13]), .B(\mem[10] [13]), .C(inst_reg[0]), 
         .Z(n37293)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32121_3_lut.init = 16'hcaca;
    LUT4 i32120_3_lut (.A(\mem[13] [13]), .B(\from_fpgacfg.wfm_ch_en [13]), 
         .C(inst_reg[0]), .Z(n37292)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32120_3_lut.init = 16'hcaca;
    LUT4 i32119_3_lut (.A(\from_fpgacfg.sync_size [13]), .B(\mem[14] [13]), 
         .C(inst_reg[0]), .Z(n37291)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32119_3_lut.init = 16'hcaca;
    LUT4 i32115_3_lut (.A(\from_fpgacfg.txant_post [13]), .B(\from_fpgacfg.txant_pre [13]), 
         .C(inst_reg[0]), .Z(n37287)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32115_3_lut.init = 16'hcaca;
    LUT4 i32114_3_lut (.A(\mem[19] [13]), .B(\mem[18] [13]), .C(inst_reg[0]), 
         .Z(n37286)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32114_3_lut.init = 16'hcaca;
    LUT4 mem_18__15__I_0_207_i7_2_lut (.A(\mem[18] [6]), .B(IO_0_c_0), .Z(\from_fpgacfg.SPI_SS [6])) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(301[35:58])
    defparam mem_18__15__I_0_207_i7_2_lut.init = 16'hbbbb;
    FD1P3DX mem_31___i11 (.D(din_reg[9]), .SP(REF_CLK_c_enable_202), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_31___i11.GSR = "ENABLED";
    FD1P3DX mem_31___i6 (.D(din_reg[4]), .SP(REF_CLK_c_enable_202), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_31___i6.GSR = "ENABLED";
    LUT4 i32113_3_lut (.A(\mem[21] [13]), .B(\mem[20] [13]), .C(inst_reg[0]), 
         .Z(n37285)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32113_3_lut.init = 16'hcaca;
    FD1P3DX mem_31___i12 (.D(din_reg[10]), .SP(REF_CLK_c_enable_202), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_31___i12.GSR = "ENABLED";
    LUT4 i32112_3_lut (.A(\from_fpgacfg.GPIO [13]), .B(\mem[22] [13]), .C(inst_reg[0]), 
         .Z(n37284)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32112_3_lut.init = 16'hcaca;
    FD1P3BX mem_31___i5 (.D(din_reg[3]), .SP(REF_CLK_c_enable_202), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.sync_pulse_period [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_31___i5.GSR = "ENABLED";
    FD1P3BX mem_31___i15 (.D(din_reg[13]), .SP(REF_CLK_c_enable_202), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.sync_pulse_period [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_31___i15.GSR = "ENABLED";
    FD1P3DX mem_30___i6 (.D(din_reg[4]), .SP(REF_CLK_c_enable_1608), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [21])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_30___i6.GSR = "ENABLED";
    FD1P3DX dout_reg_i4 (.D(dout_reg_15__N_4993[4]), .SP(sclk_N_5010_enable_16), 
            .CK(sclk_N_5010), .CD(n41434), .Q(dout_reg[4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(151[7] 170[14])
    defparam dout_reg_i4.GSR = "ENABLED";
    FD1P3DX dout_reg_i3 (.D(dout_reg_15__N_4993[3]), .SP(sclk_N_5010_enable_16), 
            .CK(sclk_N_5010), .CD(n41434), .Q(dout_reg[3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(151[7] 170[14])
    defparam dout_reg_i3.GSR = "ENABLED";
    LUT4 i32183_3_lut (.A(\mem[13] [10]), .B(\from_fpgacfg.wfm_ch_en [10]), 
         .C(inst_reg[0]), .Z(n37355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32183_3_lut.init = 16'hcaca;
    LUT4 i32182_3_lut (.A(\from_fpgacfg.sync_size [10]), .B(\mem[14] [10]), 
         .C(inst_reg[0]), .Z(n37354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32182_3_lut.init = 16'hcaca;
    FD1P3DX mem_30___i5 (.D(din_reg[3]), .SP(REF_CLK_c_enable_1608), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [20])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_30___i5.GSR = "ENABLED";
    LUT4 i32178_3_lut (.A(\from_fpgacfg.txant_post [10]), .B(\from_fpgacfg.txant_pre [10]), 
         .C(inst_reg[0]), .Z(n37350)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32178_3_lut.init = 16'hcaca;
    LUT4 i32177_3_lut (.A(\mem[19] [10]), .B(\mem[18] [10]), .C(inst_reg[0]), 
         .Z(n37349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32177_3_lut.init = 16'hcaca;
    LUT4 i32108_3_lut (.A(\mem[1] [14]), .B(\mem[0] [14]), .C(inst_reg[0]), 
         .Z(n37280)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32108_3_lut.init = 16'hcaca;
    FD1P3DX dout_reg_i2 (.D(dout_reg_15__N_4993[2]), .SP(sclk_N_5010_enable_16), 
            .CK(sclk_N_5010), .CD(n41434), .Q(dout_reg[2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(151[7] 170[14])
    defparam dout_reg_i2.GSR = "ENABLED";
    FD1P3DX dout_reg_i1 (.D(dout_reg_15__N_4993[1]), .SP(sclk_N_5010_enable_16), 
            .CK(sclk_N_5010), .CD(n41434), .Q(dout_reg[1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(151[7] 170[14])
    defparam dout_reg_i1.GSR = "ENABLED";
    FD1P3DX mem_31___i14 (.D(din_reg[12]), .SP(REF_CLK_c_enable_202), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_31___i14.GSR = "ENABLED";
    FD1P3DX mem_30___i4 (.D(din_reg[2]), .SP(REF_CLK_c_enable_1608), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [19])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_30___i4.GSR = "ENABLED";
    LUT4 i32107_3_lut (.A(\mem[3] [14]), .B(\mem[2] [14]), .C(inst_reg[0]), 
         .Z(n37279)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32107_3_lut.init = 16'hcaca;
    LUT4 i32106_3_lut (.A(\from_fpgacfg.drct_clk_en [14]), .B(\from_fpgacfg.phase_reg_sel [14]), 
         .C(inst_reg[0]), .Z(n37278)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32106_3_lut.init = 16'hcaca;
    FD1P3DX mem_30___i16 (.D(din_reg[14]), .SP(REF_CLK_c_enable_1608), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [31])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_30___i16.GSR = "ENABLED";
    LUT4 i32176_3_lut (.A(\mem[21] [10]), .B(\mem[20] [10]), .C(inst_reg[0]), 
         .Z(n37348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32176_3_lut.init = 16'hcaca;
    FD1P3DX mem_30___i15 (.D(din_reg[13]), .SP(REF_CLK_c_enable_1608), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [30])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_30___i15.GSR = "ENABLED";
    LUT4 i32175_3_lut (.A(\from_fpgacfg.GPIO [10]), .B(\mem[22] [10]), .C(inst_reg[0]), 
         .Z(n37347)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32175_3_lut.init = 16'hcaca;
    FD1P3DX mem_30___i3 (.D(din_reg[1]), .SP(REF_CLK_c_enable_1608), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [18])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_30___i3.GSR = "ENABLED";
    FD1P3DX mem_30___i14 (.D(din_reg[12]), .SP(REF_CLK_c_enable_1608), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [29])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_30___i14.GSR = "ENABLED";
    FD1P3DX mem_30___i13 (.D(din_reg[11]), .SP(REF_CLK_c_enable_1608), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [28])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_30___i13.GSR = "ENABLED";
    LUT4 i32105_3_lut (.A(\from_fpgacfg.ch_en [14]), .B(\mem[6] [14]), .C(inst_reg[0]), 
         .Z(n37277)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32105_3_lut.init = 16'hcaca;
    FD1P3DX mem_12__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_205), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.wfm_ch_en [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_12__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_12__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_205), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.wfm_ch_en [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_12__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_31___i10 (.D(din_reg[8]), .SP(REF_CLK_c_enable_202), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_31___i10.GSR = "ENABLED";
    FD1P3BX mem_12__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_205), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.wfm_ch_en [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_12__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_30___i12 (.D(din_reg[10]), .SP(REF_CLK_c_enable_1608), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [27])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_30___i12.GSR = "ENABLED";
    FD1P3DX mem_13___i16 (.D(din_reg[14]), .SP(REF_CLK_c_enable_101), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[13] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_13___i16.GSR = "ENABLED";
    FD1P3DX mem_13___i15 (.D(din_reg[13]), .SP(REF_CLK_c_enable_101), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[13] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_13___i15.GSR = "ENABLED";
    FD1P3DX mem_13___i14 (.D(din_reg[12]), .SP(REF_CLK_c_enable_101), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[13] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_13___i14.GSR = "ENABLED";
    FD1P3DX mem_13___i13 (.D(din_reg[11]), .SP(REF_CLK_c_enable_101), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[13] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_13___i13.GSR = "ENABLED";
    FD1P3BX mem_31___i13 (.D(din_reg[11]), .SP(REF_CLK_c_enable_202), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.sync_pulse_period [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_31___i13.GSR = "ENABLED";
    FD1P3DX mem_13___i12 (.D(din_reg[10]), .SP(REF_CLK_c_enable_101), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[13] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_13___i12.GSR = "ENABLED";
    FD1P3DX mem_13___i11 (.D(din_reg[9]), .SP(REF_CLK_c_enable_101), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[13] [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_13___i11.GSR = "ENABLED";
    LUT4 i32171_3_lut (.A(\mem[1] [11]), .B(\mem[0] [11]), .C(inst_reg[0]), 
         .Z(n37343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32171_3_lut.init = 16'hcaca;
    LUT4 i32170_3_lut (.A(\mem[3] [11]), .B(\mem[2] [11]), .C(inst_reg[0]), 
         .Z(n37342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32170_3_lut.init = 16'hcaca;
    LUT4 i32169_3_lut (.A(\from_fpgacfg.drct_clk_en [11]), .B(\from_fpgacfg.phase_reg_sel [11]), 
         .C(inst_reg[0]), .Z(n37341)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32169_3_lut.init = 16'hcaca;
    LUT4 i32101_3_lut (.A(\mem[9] [14]), .B(\mem[8] [14]), .C(inst_reg[0]), 
         .Z(n37273)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32101_3_lut.init = 16'hcaca;
    LUT4 i32168_3_lut (.A(\from_fpgacfg.ch_en [11]), .B(\mem[6] [11]), .C(inst_reg[0]), 
         .Z(n37340)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32168_3_lut.init = 16'hcaca;
    LUT4 i32100_3_lut (.A(\mem[11] [14]), .B(\mem[10] [14]), .C(inst_reg[0]), 
         .Z(n37272)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32100_3_lut.init = 16'hcaca;
    FD1P3DX mem_13___i10 (.D(din_reg[8]), .SP(REF_CLK_c_enable_101), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[13] [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_13___i10.GSR = "ENABLED";
    FD1P3DX mem_13___i9 (.D(din_reg[7]), .SP(REF_CLK_c_enable_101), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[13] [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_13___i9.GSR = "ENABLED";
    FD1P3DX mem_13___i8 (.D(din_reg[6]), .SP(REF_CLK_c_enable_101), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[13] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_13___i8.GSR = "ENABLED";
    LUT4 i32099_3_lut (.A(\mem[13] [14]), .B(\from_fpgacfg.wfm_ch_en [14]), 
         .C(inst_reg[0]), .Z(n37271)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32099_3_lut.init = 16'hcaca;
    LUT4 i32098_3_lut (.A(\from_fpgacfg.sync_size [14]), .B(\mem[14] [14]), 
         .C(inst_reg[0]), .Z(n37270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32098_3_lut.init = 16'hcaca;
    FD1P3DX mem_13___i7 (.D(din_reg[5]), .SP(REF_CLK_c_enable_101), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[13] [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_13___i7.GSR = "ENABLED";
    FD1P3DX mem_13___i6 (.D(din_reg[4]), .SP(REF_CLK_c_enable_101), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[13] [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_13___i6.GSR = "ENABLED";
    FD1P3BX mem_30___i2 (.D(din_reg[0]), .SP(REF_CLK_c_enable_1608), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.sync_pulse_period [17])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_30___i2.GSR = "ENABLED";
    LUT4 i15591_2_lut_rep_814 (.A(n1800[16]), .B(n11745), .Z(n41219)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i15591_2_lut_rep_814.init = 16'heeee;
    FD1P3DX mem_13___i5 (.D(din_reg[3]), .SP(REF_CLK_c_enable_101), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[13] [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_13___i5.GSR = "ENABLED";
    FD1P3DX mem_13___i4 (.D(din_reg[2]), .SP(REF_CLK_c_enable_101), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[13] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_13___i4.GSR = "ENABLED";
    FD1P3DX mem_13___i3 (.D(din_reg[1]), .SP(REF_CLK_c_enable_101), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\inst2_from_fpgacfg.wfm_load )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_13___i3.GSR = "ENABLED";
    FD1P3DX mem_13___i2 (.D(din_reg[0]), .SP(REF_CLK_c_enable_101), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\inst2_from_fpgacfg.wfm_play )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_13___i2.GSR = "ENABLED";
    FD1P3DX mem_14__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_119), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[14] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_14__i0_i15.GSR = "ENABLED";
    FD1P3DX mem_14__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_119), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[14] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_14__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_14__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_119), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[14] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_14__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_14__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_119), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[14] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_14__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_14__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_119), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[14] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_14__i0_i11.GSR = "ENABLED";
    FD1P3DX mem_14__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_119), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[14] [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_14__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_14__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_119), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[14] [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_14__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_14__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_119), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[14] [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_14__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_14__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_119), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[14] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_14__i0_i7.GSR = "ENABLED";
    FD1P3DX mem_14__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_119), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[14] [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_14__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_14__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_119), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[14] [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_14__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_14__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_119), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[14] [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_14__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_14__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_119), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[14] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_14__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_14__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_119), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[14] [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_14__i0_i2.GSR = "ENABLED";
    FD1P3BX mem_14__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_119), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[14] [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_14__i0_i1.GSR = "ENABLED";
    LUT4 i32094_3_lut (.A(\from_fpgacfg.txant_post [14]), .B(\from_fpgacfg.txant_pre [14]), 
         .C(inst_reg[0]), .Z(n37266)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32094_3_lut.init = 16'hcaca;
    FD1P3DX mem_15__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_174), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.sync_size [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_15__i0_i15.GSR = "ENABLED";
    FD1P3DX mem_30___i11 (.D(din_reg[9]), .SP(REF_CLK_c_enable_1608), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [26])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_30___i11.GSR = "ENABLED";
    LUT4 i32093_3_lut (.A(\mem[19] [14]), .B(\mem[18] [14]), .C(inst_reg[0]), 
         .Z(n37265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32093_3_lut.init = 16'hcaca;
    LUT4 i32092_3_lut (.A(\mem[21] [14]), .B(\mem[20] [14]), .C(inst_reg[0]), 
         .Z(n37264)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32092_3_lut.init = 16'hcaca;
    FD1P3DX mem_15__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_174), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.sync_size [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_15__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_30___i10 (.D(din_reg[8]), .SP(REF_CLK_c_enable_1608), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [25])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_30___i10.GSR = "ENABLED";
    FD1P3DX mem_15__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_174), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.sync_size [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_15__i0_i13.GSR = "ENABLED";
    LUT4 i32091_3_lut (.A(\from_fpgacfg.GPIO [14]), .B(\mem[22] [14]), .C(inst_reg[0]), 
         .Z(n37263)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32091_3_lut.init = 16'hcaca;
    FD1P3DX mem_15__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_174), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.sync_size [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_15__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_12__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_205), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.wfm_ch_en [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_12__i0_i15.GSR = "ENABLED";
    LUT4 i32087_3_lut (.A(\mem[1] [15]), .B(\mem[0] [15]), .C(inst_reg[0]), 
         .Z(n37259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32087_3_lut.init = 16'hcaca;
    FD1P3DX mem_31___i4 (.D(din_reg[2]), .SP(REF_CLK_c_enable_202), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_31___i4.GSR = "ENABLED";
    LUT4 i32086_3_lut (.A(\mem[3] [15]), .B(\mem[2] [15]), .C(inst_reg[0]), 
         .Z(n37258)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32086_3_lut.init = 16'hcaca;
    FD1P3BX mem_31___i16 (.D(din_reg[14]), .SP(REF_CLK_c_enable_202), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.sync_pulse_period [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_31___i16.GSR = "ENABLED";
    FD1P3DX mem_15__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_174), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.sync_size [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_15__i0_i11.GSR = "ENABLED";
    LUT4 i32085_3_lut (.A(\from_fpgacfg.drct_clk_en [15]), .B(\from_fpgacfg.phase_reg_sel [15]), 
         .C(inst_reg[0]), .Z(n37257)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32085_3_lut.init = 16'hcaca;
    FD1P3DX mem_30___i9 (.D(din_reg[7]), .SP(REF_CLK_c_enable_1608), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [24])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_30___i9.GSR = "ENABLED";
    FD1P3DX mem_15__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_174), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_size [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_15__i0_i10.GSR = "ENABLED";
    FD1P3BX mem_15__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_174), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.sync_size [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_15__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_30___i8 (.D(din_reg[6]), .SP(REF_CLK_c_enable_1608), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [23])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_30___i8.GSR = "ENABLED";
    LUT4 i32084_3_lut (.A(\from_fpgacfg.ch_en [15]), .B(\mem[6] [15]), .C(inst_reg[0]), 
         .Z(n37256)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32084_3_lut.init = 16'hcaca;
    LUT4 i32080_3_lut (.A(\mem[9] [15]), .B(\mem[8] [15]), .C(inst_reg[0]), 
         .Z(n37252)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32080_3_lut.init = 16'hcaca;
    FD1P3BX mem_15__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_174), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.sync_size [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_15__i0_i8.GSR = "ENABLED";
    LUT4 i32164_3_lut (.A(\mem[9] [11]), .B(\mem[8] [11]), .C(inst_reg[0]), 
         .Z(n37336)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32164_3_lut.init = 16'hcaca;
    FD1P3DX mem_12__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_205), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.wfm_ch_en [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_12__i0_i14.GSR = "ENABLED";
    LUT4 i32079_3_lut (.A(\mem[11] [15]), .B(\mem[10] [15]), .C(inst_reg[0]), 
         .Z(n37251)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32079_3_lut.init = 16'hcaca;
    LUT4 i32078_3_lut (.A(\mem[13] [15]), .B(\from_fpgacfg.wfm_ch_en [15]), 
         .C(inst_reg[0]), .Z(n37250)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32078_3_lut.init = 16'hcaca;
    FD1P3BX mem_15__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_174), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.sync_size [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_15__i0_i7.GSR = "ENABLED";
    LUT4 i32163_3_lut (.A(\mem[11] [11]), .B(\mem[10] [11]), .C(inst_reg[0]), 
         .Z(n37335)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32163_3_lut.init = 16'hcaca;
    FD1P3BX mem_15__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_174), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.sync_size [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_15__i0_i6.GSR = "ENABLED";
    LUT4 mux_16_Mux_2_i27_3_lut (.A(\mem[1] [2]), .B(\mem[0] [2]), .C(inst_reg[0]), 
         .Z(n27)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam mux_16_Mux_2_i27_3_lut.init = 16'hcaca;
    FD1P3BX mem_15__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_174), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.sync_size [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_15__i0_i5.GSR = "ENABLED";
    FD1P3BX mem_15__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_174), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.sync_size [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_15__i0_i4.GSR = "ENABLED";
    FD1P3BX mem_15__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_174), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.sync_size [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_15__i0_i3.GSR = "ENABLED";
    FD1P3BX mem_15__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_174), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.sync_size [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_15__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_15__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_174), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_size [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_15__i0_i1.GSR = "ENABLED";
    LUT4 mem_18__15__I_0_207_i6_2_lut (.A(\mem[18] [5]), .B(IO_0_c_0), .Z(\from_fpgacfg.SPI_SS [5])) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(301[35:58])
    defparam mem_18__15__I_0_207_i6_2_lut.init = 16'hbbbb;
    FD1P3DX mem_16__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_211), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.txant_pre [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_16__i0_i15.GSR = "ENABLED";
    FD1P3DX inst_reg_i0_i0 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_1424), .CK(REF_CLK_c), 
            .CD(n41434), .Q(inst_reg[0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(115[7] 124[14])
    defparam inst_reg_i0_i0.GSR = "ENABLED";
    FD1P3DX mem_16__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_211), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.txant_pre [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_16__i0_i14.GSR = "ENABLED";
    LUT4 i32077_3_lut (.A(\from_fpgacfg.sync_size [15]), .B(\mem[14] [15]), 
         .C(inst_reg[0]), .Z(n37249)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32077_3_lut.init = 16'hcaca;
    FD1P3DX mem_16__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_211), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.txant_pre [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_16__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_16__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_211), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.txant_pre [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_16__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_12__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_205), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.wfm_ch_en [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_12__i0_i13.GSR = "ENABLED";
    LUT4 mem_18__15__I_0_207_i5_2_lut (.A(\mem[18] [4]), .B(IO_0_c_0), .Z(\from_fpgacfg.SPI_SS [4])) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(301[35:58])
    defparam mem_18__15__I_0_207_i5_2_lut.init = 16'hbbbb;
    FD1P3DX mem_16__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_211), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.txant_pre [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_16__i0_i11.GSR = "ENABLED";
    LUT4 i32073_3_lut (.A(\from_fpgacfg.txant_post [15]), .B(\from_fpgacfg.txant_pre [15]), 
         .C(inst_reg[0]), .Z(n37245)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32073_3_lut.init = 16'hcaca;
    FD1P3DX mem_16__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_211), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_pre [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_16__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_31___i9 (.D(din_reg[7]), .SP(REF_CLK_c_enable_202), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_31___i9.GSR = "ENABLED";
    LUT4 i32162_3_lut (.A(\mem[13] [11]), .B(\from_fpgacfg.wfm_ch_en [11]), 
         .C(inst_reg[0]), .Z(n37334)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32162_3_lut.init = 16'hcaca;
    LUT4 i32161_3_lut (.A(\from_fpgacfg.sync_size [11]), .B(\mem[14] [11]), 
         .C(inst_reg[0]), .Z(n37333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32161_3_lut.init = 16'hcaca;
    LUT4 i32072_3_lut (.A(\mem[19] [15]), .B(\mem[18] [15]), .C(inst_reg[0]), 
         .Z(n37244)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32072_3_lut.init = 16'hcaca;
    LUT4 i32157_3_lut (.A(\from_fpgacfg.txant_post [11]), .B(\from_fpgacfg.txant_pre [11]), 
         .C(inst_reg[0]), .Z(n37329)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32157_3_lut.init = 16'hcaca;
    LUT4 i32156_3_lut (.A(\mem[19] [11]), .B(\mem[18] [11]), .C(inst_reg[0]), 
         .Z(n37328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32156_3_lut.init = 16'hcaca;
    FD1P3DX mem_31___i3 (.D(din_reg[1]), .SP(REF_CLK_c_enable_202), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_31___i3.GSR = "ENABLED";
    LUT4 i32071_3_lut (.A(\mem[21] [15]), .B(\mem[20] [15]), .C(inst_reg[0]), 
         .Z(n37243)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32071_3_lut.init = 16'hcaca;
    FD1P3DX mem_31___i2 (.D(din_reg[0]), .SP(REF_CLK_c_enable_202), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_31___i2.GSR = "ENABLED";
    FD1P3DX mem_31___i1 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_202), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_31___i1.GSR = "ENABLED";
    LUT4 i32070_3_lut (.A(\from_fpgacfg.GPIO [15]), .B(\mem[22] [15]), .C(inst_reg[0]), 
         .Z(n37242)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32070_3_lut.init = 16'hcaca;
    LUT4 i32155_3_lut (.A(\mem[21] [11]), .B(\mem[20] [11]), .C(inst_reg[0]), 
         .Z(n37327)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32155_3_lut.init = 16'hcaca;
    FD1P3DX mem_16__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_211), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_pre [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_16__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_16__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_211), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_pre [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_16__i0_i8.GSR = "ENABLED";
    LUT4 i32154_3_lut (.A(\from_fpgacfg.GPIO [11]), .B(\mem[22] [11]), .C(inst_reg[0]), 
         .Z(n37326)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32154_3_lut.init = 16'hcaca;
    FD1P3DX mem_16__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_211), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_pre [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_16__i0_i7.GSR = "ENABLED";
    LUT4 i32150_3_lut (.A(\mem[1] [12]), .B(\mem[0] [12]), .C(inst_reg[0]), 
         .Z(n37322)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32150_3_lut.init = 16'hcaca;
    FD1P3BX mem_31___i8 (.D(din_reg[6]), .SP(REF_CLK_c_enable_202), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.sync_pulse_period [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_31___i8.GSR = "ENABLED";
    FD1P3DX mem_16__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_211), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_pre [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_16__i0_i6.GSR = "ENABLED";
    LUT4 i32149_3_lut (.A(\mem[3] [12]), .B(\mem[2] [12]), .C(inst_reg[0]), 
         .Z(n37321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32149_3_lut.init = 16'hcaca;
    LUT4 mem_18__15__I_0_207_i10_2_lut (.A(\mem[18] [9]), .B(IO_0_c_0), 
         .Z(\from_fpgacfg.SPI_SS [9])) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(301[35:58])
    defparam mem_18__15__I_0_207_i10_2_lut.init = 16'hbbbb;
    LUT4 i32148_3_lut (.A(\from_fpgacfg.drct_clk_en [12]), .B(\from_fpgacfg.phase_reg_sel [12]), 
         .C(inst_reg[0]), .Z(n37320)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32148_3_lut.init = 16'hcaca;
    LUT4 i32147_3_lut (.A(\from_fpgacfg.ch_en [12]), .B(\mem[6] [12]), .C(inst_reg[0]), 
         .Z(n37319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32147_3_lut.init = 16'hcaca;
    FD1P3DX mem_31___i7 (.D(din_reg[5]), .SP(REF_CLK_c_enable_202), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_31___i7.GSR = "ENABLED";
    PFUMX i34357 (.BLUT(n41456), .ALUT(n41457), .C0(inst_reg[0]), .Z(n41458));
    FD1P3DX mem_16__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_211), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_pre [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_16__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_12__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_205), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.wfm_ch_en [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_12__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_12__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_205), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.wfm_ch_en [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_12__i0_i11.GSR = "ENABLED";
    LUT4 mem_18__15__I_0_207_i4_2_lut (.A(\mem[18] [3]), .B(IO_0_c_0), .Z(\from_fpgacfg.SPI_SS [3])) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(301[35:58])
    defparam mem_18__15__I_0_207_i4_2_lut.init = 16'hbbbb;
    FD1P3DX mem_16__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_211), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_pre [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_16__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_16__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_211), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_pre [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_16__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_16__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_211), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_pre [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_16__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_16__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_211), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_pre [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_16__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_17__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_226), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.txant_post [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_17__i0_i15.GSR = "ENABLED";
    FD1P3DX mem_17__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_226), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.txant_post [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_17__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_17__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_226), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.txant_post [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_17__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_17__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_226), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.txant_post [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_17__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_17__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_226), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.txant_post [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_17__i0_i11.GSR = "ENABLED";
    FD1P3DX mem_17__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_226), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_post [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_17__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_17__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_226), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_post [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_17__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_17__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_226), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_post [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_17__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_17__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_226), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_post [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_17__i0_i7.GSR = "ENABLED";
    FD1P3DX mem_17__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_226), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_post [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_17__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_17__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_226), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_post [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_17__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_17__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_226), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_post [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_17__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_17__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_226), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_post [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_17__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_17__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_226), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_post [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_17__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_17__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_226), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.txant_post [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_17__i0_i1.GSR = "ENABLED";
    FD1P3BX mem_18__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_242), 
            .CK(REF_CLK_c), .PD(n41434), .Q(\mem[18] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_18__i0_i15.GSR = "ENABLED";
    FD1P3BX mem_18__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_242), 
            .CK(REF_CLK_c), .PD(n41434), .Q(\mem[18] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_18__i0_i14.GSR = "ENABLED";
    FD1P3BX mem_18__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_242), 
            .CK(REF_CLK_c), .PD(n41434), .Q(\mem[18] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_18__i0_i13.GSR = "ENABLED";
    FD1P3BX mem_18__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_242), 
            .CK(REF_CLK_c), .PD(n41434), .Q(\mem[18] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_18__i0_i12.GSR = "ENABLED";
    FD1P3BX mem_18__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_242), 
            .CK(REF_CLK_c), .PD(n41434), .Q(\mem[18] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_18__i0_i11.GSR = "ENABLED";
    FD1P3BX mem_18__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_242), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[18] [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_18__i0_i10.GSR = "ENABLED";
    FD1P3BX mem_18__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_242), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[18] [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_18__i0_i9.GSR = "ENABLED";
    FD1P3BX mem_18__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_242), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[18] [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_18__i0_i8.GSR = "ENABLED";
    FD1P3BX mem_18__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_242), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[18] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_18__i0_i7.GSR = "ENABLED";
    FD1P3BX mem_18__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_242), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[18] [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_18__i0_i6.GSR = "ENABLED";
    FD1P3BX mem_18__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_242), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[18] [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_18__i0_i5.GSR = "ENABLED";
    FD1P3BX mem_18__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_242), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[18] [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_18__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_30___i7 (.D(din_reg[5]), .SP(REF_CLK_c_enable_1608), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.sync_pulse_period [22])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_30___i7.GSR = "ENABLED";
    FD1P3BX mem_18__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_242), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[18] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_18__i0_i3.GSR = "ENABLED";
    FD1P3BX mem_18__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_242), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[18] [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_18__i0_i2.GSR = "ENABLED";
    FD1P3BX mem_18__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_242), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[18] [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_18__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_19__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_258), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[19] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_19__i0_i15.GSR = "ENABLED";
    FD1P3BX mem_19__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_258), 
            .CK(REF_CLK_c), .PD(n41434), .Q(\mem[19] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_19__i0_i14.GSR = "ENABLED";
    FD1P3BX mem_19__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_258), 
            .CK(REF_CLK_c), .PD(n41434), .Q(\mem[19] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_19__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_19__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_258), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[19] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_19__i0_i12.GSR = "ENABLED";
    FD1P3BX mem_19__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_258), 
            .CK(REF_CLK_c), .PD(n41434), .Q(\mem[19] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_19__i0_i11.GSR = "ENABLED";
    FD1P3BX mem_19__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_258), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[19] [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_19__i0_i10.GSR = "ENABLED";
    FD1P3BX mem_19__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_258), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[19] [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_19__i0_i9.GSR = "ENABLED";
    FD1P3BX mem_19__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_258), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[19] [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_19__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_19__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_258), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[19] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_19__i0_i7.GSR = "ENABLED";
    FD1P3BX mem_19__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_258), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\inst2_from_fpgacfg.LMS1_RXEN )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_19__i0_i6.GSR = "ENABLED";
    FD1P3BX mem_19__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_258), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\inst2_from_fpgacfg.LMS1_TXEN )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_19__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_19__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_258), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\inst2_from_fpgacfg.LMS1_TXNRX2 )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_19__i0_i4.GSR = "ENABLED";
    FD1P3BX mem_19__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_258), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\inst2_from_fpgacfg.LMS1_TXNRX1 )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_19__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_19__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_258), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\inst2_from_fpgacfg.LMS1_CORE_LDO_EN )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_19__i0_i2.GSR = "ENABLED";
    FD1P3BX mem_19__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_258), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\inst2_from_fpgacfg.LMS1_RESET )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_19__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_20__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_273), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[20] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_20__i0_i15.GSR = "ENABLED";
    FD1P3DX mem_20__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_273), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[20] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_20__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_20__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_273), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[20] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_20__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_20__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_273), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[20] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_20__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_20__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_273), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[20] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_20__i0_i11.GSR = "ENABLED";
    FD1P3DX mem_20__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_273), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[20] [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_20__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_20__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_273), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[20] [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_20__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_20__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_273), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[20] [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_20__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_20__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_273), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[20] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_20__i0_i7.GSR = "ENABLED";
    FD1P3DX mem_20__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_273), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[20] [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_20__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_20__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_273), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[20] [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_20__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_20__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_273), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[20] [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_20__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_20__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_273), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[20] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_20__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_20__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_273), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[20] [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_20__i0_i2.GSR = "ENABLED";
    FD1P3BX mem_20__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_273), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\mem[20] [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_20__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_21__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_289), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[21] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_21__i0_i15.GSR = "ENABLED";
    FD1P3DX mem_21__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_289), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[21] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_21__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_21__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_289), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[21] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_21__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_21__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_289), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[21] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_21__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_21__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_289), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[21] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_21__i0_i11.GSR = "ENABLED";
    FD1P3DX mem_21__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_289), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[21] [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_21__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_21__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_289), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[21] [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_21__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_21__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_289), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[21] [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_21__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_21__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_289), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[21] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_21__i0_i7.GSR = "ENABLED";
    LUT4 mem_18__15__I_0_207_i3_2_lut (.A(\mem[18] [2]), .B(IO_0_c_0), .Z(\from_fpgacfg.SPI_SS [2])) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(301[35:58])
    defparam mem_18__15__I_0_207_i3_2_lut.init = 16'hbbbb;
    FD1P3DX mem_21__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_289), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[21] [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_21__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_21__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_289), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[21] [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_21__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_21__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_289), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[21] [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_21__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_21__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_289), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[21] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_21__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_21__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_289), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[21] [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_21__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_21__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_289), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[21] [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_21__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_22__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_304), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[22] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_22__i0_i15.GSR = "ENABLED";
    FD1P3DX mem_22__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_304), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[22] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_22__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_22__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_304), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[22] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_22__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_22__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_304), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[22] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_22__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_22__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_304), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[22] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_22__i0_i11.GSR = "ENABLED";
    FD1P3DX mem_22__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_304), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[22] [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_22__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_22__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_304), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[22] [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_22__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_22__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_304), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[22] [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_22__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_22__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_304), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[22] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_22__i0_i7.GSR = "ENABLED";
    FD1P3DX mem_22__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_304), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[22] [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_22__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_22__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_304), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[22] [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_22__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_22__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_304), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[22] [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_22__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_22__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_304), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[22] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_22__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_22__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_304), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[22] [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_22__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_22__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_304), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[22] [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_22__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_23__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_322), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.GPIO [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_23__i0_i15.GSR = "ENABLED";
    FD1P3DX mem_23__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_322), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.GPIO [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_23__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_23__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_322), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.GPIO [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_23__i0_i13.GSR = "ENABLED";
    FD1P3BX mem_23__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_322), 
            .CK(REF_CLK_c), .PD(n41434), .Q(\from_fpgacfg.GPIO [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_23__i0_i12.GSR = "ENABLED";
    LUT4 i31142_3_lut (.A(\mem[25] [12]), .B(\mem[24] [12]), .C(inst_reg[0]), 
         .Z(n36314)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31142_3_lut.init = 16'hcaca;
    FD1P3DX mem_23__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_322), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\from_fpgacfg.GPIO [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_23__i0_i11.GSR = "ENABLED";
    LUT4 i31141_3_lut (.A(\mem[27] [12]), .B(\mem[26] [12]), .C(inst_reg[0]), 
         .Z(n36313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31141_3_lut.init = 16'hcaca;
    FD1P3DX mem_23__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_322), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.GPIO [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_23__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_23__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_322), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.GPIO [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_23__i0_i9.GSR = "ENABLED";
    FD1P3BX mem_23__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_322), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.GPIO [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_23__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_23__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_322), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.GPIO [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_23__i0_i7.GSR = "ENABLED";
    FD1P3BX mem_23__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_322), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.GPIO [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_23__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_23__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_322), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.GPIO [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_23__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_23__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_322), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.GPIO [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_23__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_23__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_322), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.GPIO [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_23__i0_i3.GSR = "ENABLED";
    FD1P3BX mem_23__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_322), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.GPIO [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_23__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_23__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_322), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.GPIO [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_23__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_24__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_337), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[24] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_24__i0_i15.GSR = "ENABLED";
    FD1P3DX mem_24__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_337), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[24] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_24__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_24__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_337), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[24] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_24__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_24__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_337), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[24] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_24__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_24__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_337), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[24] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_24__i0_i11.GSR = "ENABLED";
    FD1P3DX mem_24__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_337), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[24] [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_24__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_24__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_337), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[24] [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_24__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_24__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_337), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[24] [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_24__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_24__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_337), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[24] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_24__i0_i7.GSR = "ENABLED";
    FD1P3DX mem_24__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_337), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[24] [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_24__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_24__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_337), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[24] [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_24__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_24__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_337), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[24] [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_24__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_24__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_337), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[24] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_24__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_24__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_337), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[24] [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_24__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_24__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_337), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[24] [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_24__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_25__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_352), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[25] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_25__i0_i15.GSR = "ENABLED";
    FD1P3DX mem_25__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_352), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[25] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_25__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_25__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_352), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[25] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_25__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_25__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_352), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[25] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_25__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_25__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_352), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[25] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_25__i0_i11.GSR = "ENABLED";
    LUT4 mem_18__15__I_0_207_i2_2_lut (.A(\mem[18] [1]), .B(IO_0_c_0), .Z(\from_fpgacfg.SPI_SS [1])) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(301[35:58])
    defparam mem_18__15__I_0_207_i2_2_lut.init = 16'hbbbb;
    PFUMX i34355 (.BLUT(n41453), .ALUT(n41454), .C0(inst_reg[0]), .Z(n41455));
    FD1P3DX mem_25__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_352), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[25] [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_25__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_25__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_352), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[25] [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_25__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_25__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_352), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[25] [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_25__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_25__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_352), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[25] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_25__i0_i7.GSR = "ENABLED";
    FD1P3DX mem_25__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_352), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[25] [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_25__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_25__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_352), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[25] [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_25__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_25__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_352), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[25] [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_25__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_25__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_352), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[25] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_25__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_25__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_352), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[25] [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_25__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_25__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_352), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[25] [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_25__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_26___i16 (.D(din_reg[14]), .SP(REF_CLK_c_enable_367), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[26] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_26___i16.GSR = "ENABLED";
    FD1P3DX mem_26___i15 (.D(din_reg[13]), .SP(REF_CLK_c_enable_367), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[26] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_26___i15.GSR = "ENABLED";
    FD1P3DX mem_26___i14 (.D(din_reg[12]), .SP(REF_CLK_c_enable_367), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[26] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_26___i14.GSR = "ENABLED";
    FD1P3DX mem_26___i13 (.D(din_reg[11]), .SP(REF_CLK_c_enable_367), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[26] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_26___i13.GSR = "ENABLED";
    FD1P3DX mem_26___i12 (.D(din_reg[10]), .SP(REF_CLK_c_enable_367), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[26] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_26___i12.GSR = "ENABLED";
    FD1P3DX mem_26___i11 (.D(din_reg[9]), .SP(REF_CLK_c_enable_367), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[26] [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_26___i11.GSR = "ENABLED";
    FD1P3DX mem_26___i10 (.D(din_reg[8]), .SP(REF_CLK_c_enable_367), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[26] [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_26___i10.GSR = "ENABLED";
    FD1P3DX mem_26___i9 (.D(din_reg[7]), .SP(REF_CLK_c_enable_367), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[26] [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_26___i9.GSR = "ENABLED";
    FD1P3DX mem_26___i8 (.D(din_reg[6]), .SP(REF_CLK_c_enable_367), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[26] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_26___i8.GSR = "ENABLED";
    FD1P3DX mem_26___i7 (.D(din_reg[5]), .SP(REF_CLK_c_enable_367), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.FPGA_LED2_CTRL [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_26___i7.GSR = "ENABLED";
    FD1P3DX mem_26___i6 (.D(din_reg[4]), .SP(REF_CLK_c_enable_367), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.FPGA_LED2_CTRL [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_26___i6.GSR = "ENABLED";
    FD1P3DX mem_26___i5 (.D(din_reg[3]), .SP(REF_CLK_c_enable_367), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.FPGA_LED2_CTRL [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_26___i5.GSR = "ENABLED";
    FD1P3DX mem_26___i4 (.D(din_reg[2]), .SP(REF_CLK_c_enable_367), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[26] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_26___i4.GSR = "ENABLED";
    FD1P3DX mem_26___i3 (.D(din_reg[1]), .SP(REF_CLK_c_enable_367), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.FPGA_LED1_CTRL [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_26___i3.GSR = "ENABLED";
    FD1P3DX mem_26___i2 (.D(din_reg[0]), .SP(REF_CLK_c_enable_367), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.FPGA_LED1_CTRL [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_26___i2.GSR = "ENABLED";
    FD1P3DX mem_27__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_382), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[27] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_27__i0_i15.GSR = "ENABLED";
    FD1P3DX mem_27__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_382), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[27] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_27__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_27__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_382), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[27] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_27__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_27__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_382), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[27] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_27__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_27__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_382), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[27] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_27__i0_i11.GSR = "ENABLED";
    FD1P3DX mem_27__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_382), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[27] [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_27__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_27__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_382), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[27] [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_27__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_27__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_382), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[27] [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_27__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_27__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_382), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[27] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_27__i0_i7.GSR = "ENABLED";
    FD1P3DX mem_27__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_382), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[27] [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_27__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_27__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_382), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[27] [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_27__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_27__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_382), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[27] [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_27__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_27__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_382), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[27] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_27__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_27__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_382), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[27] [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_27__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_27__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_382), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[27] [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_27__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_28__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_384), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.FX3_LED_CTRL [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_28__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_28__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_384), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.FX3_LED_CTRL [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_28__i0_i1.GSR = "ENABLED";
    FD1P3BX mem_29__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_387), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.CLK_ENA [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_29__i0_i3.GSR = "ENABLED";
    FD1P3BX mem_29__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_387), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.CLK_ENA [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_29__i0_i2.GSR = "ENABLED";
    FD1P3BX mem_29__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_387), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.CLK_ENA [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_29__i0_i1.GSR = "ENABLED";
    L6MUX21 i30785 (.D0(n37318), .D1(n37325), .SD(inst_reg[3]), .Z(n35957));
    L6MUX21 i30839 (.D0(n37339), .D1(n37346), .SD(inst_reg[3]), .Z(n36011));
    L6MUX21 i30854 (.D0(n37360), .D1(n37367), .SD(inst_reg[3]), .Z(n36026));
    LUT4 mem_18__15__I_0_207_i1_2_lut (.A(\mem[18] [0]), .B(IO_0_c_0), .Z(\from_fpgacfg.SPI_SS [0])) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(301[35:58])
    defparam mem_18__15__I_0_207_i1_2_lut.init = 16'hbbbb;
    L6MUX21 i31103 (.D0(n37255), .D1(n37262), .SD(inst_reg[3]), .Z(n36275));
    L6MUX21 i31115 (.D0(n37381), .D1(n37388), .SD(inst_reg[3]), .Z(n36287));
    L6MUX21 i31118 (.D0(n37402), .D1(n37409), .SD(inst_reg[3]), .Z(n36290));
    L6MUX21 i32024 (.D0(n37193), .D1(n37194), .SD(inst_reg[3]), .Z(n37196));
    LUT4 mem_19__0__I_0_2_lut (.A(\mem[19] [0]), .B(IO_0_c_0), .Z(\inst2_from_fpgacfg.LMS1_SS )) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(304[43:66])
    defparam mem_19__0__I_0_2_lut.init = 16'hbbbb;
    L6MUX21 i30878 (.D0(n37465), .D1(n37472), .SD(inst_reg[3]), .Z(n36050));
    L6MUX21 i32031 (.D0(n37200), .D1(n37201), .SD(inst_reg[3]), .Z(n37203));
    L6MUX21 i31124 (.D0(n37423), .D1(n37430), .SD(inst_reg[3]), .Z(n36296));
    L6MUX21 i31127 (.D0(n37444), .D1(n37451), .SD(inst_reg[3]), .Z(n36299));
    L6MUX21 i32038 (.D0(n37207), .D1(n37208), .SD(inst_reg[3]), .Z(n37210));
    L6MUX21 i31130 (.D0(n37276), .D1(n37283), .SD(inst_reg[3]), .Z(n36302));
    L6MUX21 i31139 (.D0(n37297), .D1(n37304), .SD(inst_reg[3]), .Z(n36311));
    L6MUX21 i32314 (.D0(n37483), .D1(n37484), .SD(inst_reg[3]), .Z(n37486));
    L6MUX21 i32321 (.D0(n37490), .D1(n37491), .SD(inst_reg[3]), .Z(n37493));
    L6MUX21 i32020 (.D0(n35985), .D1(n35988), .SD(inst_reg[2]), .Z(n37192));
    L6MUX21 i32021 (.D0(n35991), .D1(n35994), .SD(inst_reg[2]), .Z(n37193));
    L6MUX21 i32022 (.D0(n35997), .D1(n36000), .SD(inst_reg[2]), .Z(n37194));
    L6MUX21 i32027 (.D0(n36006), .D1(n36009), .SD(inst_reg[2]), .Z(n37199));
    L6MUX21 i32028 (.D0(n36015), .D1(n36018), .SD(inst_reg[2]), .Z(n37200));
    L6MUX21 i32029 (.D0(n36021), .D1(n36024), .SD(inst_reg[2]), .Z(n37201));
    L6MUX21 i32034 (.D0(n36033), .D1(n36036), .SD(inst_reg[2]), .Z(n37206));
    FD1P3DX din_reg__i1 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_1621), .CK(REF_CLK_c), 
            .CD(n41434), .Q(din_reg[0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(133[7] 142[14])
    defparam din_reg__i1.GSR = "ENABLED";
    L6MUX21 i32035 (.D0(n36039), .D1(n36042), .SD(inst_reg[2]), .Z(n37207));
    L6MUX21 i32036 (.D0(n36045), .D1(n36048), .SD(inst_reg[2]), .Z(n37208));
    L6MUX21 i32076 (.D0(n37246), .D1(n37247), .SD(inst_reg[2]), .Z(n37248));
    L6MUX21 i32083 (.D0(n37253), .D1(n37254), .SD(inst_reg[2]), .Z(n37255));
    L6MUX21 i32090 (.D0(n37260), .D1(n37261), .SD(inst_reg[2]), .Z(n37262));
    L6MUX21 i32097 (.D0(n37267), .D1(n37268), .SD(inst_reg[2]), .Z(n37269));
    L6MUX21 i32104 (.D0(n37274), .D1(n37275), .SD(inst_reg[2]), .Z(n37276));
    L6MUX21 i32111 (.D0(n37281), .D1(n37282), .SD(inst_reg[2]), .Z(n37283));
    L6MUX21 i32118 (.D0(n37288), .D1(n37289), .SD(inst_reg[2]), .Z(n37290));
    L6MUX21 i32125 (.D0(n37295), .D1(n37296), .SD(inst_reg[2]), .Z(n37297));
    L6MUX21 i32132 (.D0(n37302), .D1(n37303), .SD(inst_reg[2]), .Z(n37304));
    L6MUX21 i32139 (.D0(n37309), .D1(n37310), .SD(inst_reg[2]), .Z(n37311));
    FD1P3DX mem_11__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_511), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[11] [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_11__i0_i1.GSR = "ENABLED";
    FD1P3DX dout_reg_i15 (.D(dout_reg_15__N_4993[15]), .SP(sclk_N_5010_enable_16), 
            .CK(sclk_N_5010), .CD(n41434), .Q(dout_reg[15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(151[7] 170[14])
    defparam dout_reg_i15.GSR = "ENABLED";
    L6MUX21 i32146 (.D0(n37316), .D1(n37317), .SD(inst_reg[2]), .Z(n37318));
    FD1P3DX dout_reg_i14 (.D(dout_reg_15__N_4993[14]), .SP(sclk_N_5010_enable_16), 
            .CK(sclk_N_5010), .CD(n41434), .Q(dout_reg[14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(151[7] 170[14])
    defparam dout_reg_i14.GSR = "ENABLED";
    FD1P3DX dout_reg_i13 (.D(dout_reg_15__N_4993[13]), .SP(sclk_N_5010_enable_16), 
            .CK(sclk_N_5010), .CD(n41434), .Q(dout_reg[13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(151[7] 170[14])
    defparam dout_reg_i13.GSR = "ENABLED";
    FD1P3DX dout_reg_i12 (.D(dout_reg_15__N_4993[12]), .SP(sclk_N_5010_enable_16), 
            .CK(sclk_N_5010), .CD(n41434), .Q(dout_reg[12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(151[7] 170[14])
    defparam dout_reg_i12.GSR = "ENABLED";
    FD1P3DX dout_reg_i11 (.D(dout_reg_15__N_4993[11]), .SP(sclk_N_5010_enable_16), 
            .CK(sclk_N_5010), .CD(n41434), .Q(dout_reg[11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(151[7] 170[14])
    defparam dout_reg_i11.GSR = "ENABLED";
    FD1P3DX dout_reg_i10 (.D(dout_reg_15__N_4993[10]), .SP(sclk_N_5010_enable_16), 
            .CK(sclk_N_5010), .CD(n41434), .Q(dout_reg[10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(151[7] 170[14])
    defparam dout_reg_i10.GSR = "ENABLED";
    FD1P3DX dout_reg_i9 (.D(dout_reg_15__N_4993[9]), .SP(sclk_N_5010_enable_16), 
            .CK(sclk_N_5010), .CD(n41434), .Q(dout_reg[9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(151[7] 170[14])
    defparam dout_reg_i9.GSR = "ENABLED";
    FD1P3DX dout_reg_i8 (.D(dout_reg_15__N_4993[8]), .SP(sclk_N_5010_enable_16), 
            .CK(sclk_N_5010), .CD(n41434), .Q(dout_reg[8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(151[7] 170[14])
    defparam dout_reg_i8.GSR = "ENABLED";
    FD1P3DX dout_reg_i7 (.D(dout_reg_15__N_4993[7]), .SP(sclk_N_5010_enable_16), 
            .CK(sclk_N_5010), .CD(n41434), .Q(dout_reg[7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(151[7] 170[14])
    defparam dout_reg_i7.GSR = "ENABLED";
    FD1P3DX dout_reg_i6 (.D(dout_reg_15__N_4993[6]), .SP(sclk_N_5010_enable_16), 
            .CK(sclk_N_5010), .CD(n41434), .Q(dout_reg[6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(151[7] 170[14])
    defparam dout_reg_i6.GSR = "ENABLED";
    FD1P3DX dout_reg_i5 (.D(dout_reg_15__N_4993[5]), .SP(sclk_N_5010_enable_16), 
            .CK(sclk_N_5010), .CD(n41434), .Q(dout_reg[5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(151[7] 170[14])
    defparam dout_reg_i5.GSR = "ENABLED";
    FD1P3DX mem_11__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_511), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[11] [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_11__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_11__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_511), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[11] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_11__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_11__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_511), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[11] [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_11__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_11__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_511), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[11] [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_11__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_11__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_511), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[11] [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_11__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_11__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_511), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[11] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_11__i0_i7.GSR = "ENABLED";
    FD1P3DX mem_11__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_511), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[11] [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_11__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_11__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_511), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[11] [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_11__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_11__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_511), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[11] [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_11__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_11__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_511), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[11] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_11__i0_i11.GSR = "ENABLED";
    FD1P3DX mem_11__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_511), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[11] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_11__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_11__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_511), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[11] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_11__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_11__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_511), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[11] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_11__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_11__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_511), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\mem[11] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_11__i0_i15.GSR = "ENABLED";
    FD1P3DX mem_10___i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_526), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\inst2_from_fpgacfg.tx_en )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_10___i1.GSR = "ENABLED";
    FD1P3DX mem_10___i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_526), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[10] [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_10___i2.GSR = "ENABLED";
    FD1P3DX mem_10___i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_526), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[10] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_10___i3.GSR = "ENABLED";
    FD1P3DX mem_10___i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_526), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[10] [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_10___i4.GSR = "ENABLED";
    FD1P3DX mem_10___i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_526), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[10] [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_10___i5.GSR = "ENABLED";
    FD1P3DX mem_10___i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_526), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[10] [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_10___i6.GSR = "ENABLED";
    FD1P3DX mem_10___i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_526), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[10] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_10___i7.GSR = "ENABLED";
    FD1P3DX mem_10___i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_526), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\inst2_from_fpgacfg.rx_ptrn_en )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_10___i8.GSR = "ENABLED";
    FD1P3DX mem_10___i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_526), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\inst2_from_fpgacfg.tx_ptrn_en )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_10___i9.GSR = "ENABLED";
    FD1P3DX mem_10___i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_526), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\inst2_from_fpgacfg.tx_cnt_en )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_10___i10.GSR = "ENABLED";
    FD1P3DX mem_10___i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_526), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[10] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_10___i11.GSR = "ENABLED";
    FD1P3DX mem_10___i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_526), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[10] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_10___i12.GSR = "ENABLED";
    FD1P3DX mem_10___i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_526), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[10] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_10___i13.GSR = "ENABLED";
    FD1P3DX mem_10___i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_526), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[10] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_10___i14.GSR = "ENABLED";
    FD1P3DX mem_10___i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_526), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[10] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_10___i15.GSR = "ENABLED";
    FD1P3BX mem_9___i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_541), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\inst2_from_fpgacfg.txpct_loss_clr )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_9___i1.GSR = "ENABLED";
    FD1P3DX mem_9___i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_541), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[9] [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_9___i2.GSR = "ENABLED";
    FD1P3DX mem_9___i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_541), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[9] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_9___i3.GSR = "ENABLED";
    FD1P3DX mem_9___i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_541), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[9] [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_9___i4.GSR = "ENABLED";
    FD1P3DX mem_9___i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_541), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[9] [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_9___i5.GSR = "ENABLED";
    FD1P3DX mem_9___i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_541), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[9] [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_9___i6.GSR = "ENABLED";
    FD1P3DX mem_9___i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_541), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[9] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_9___i7.GSR = "ENABLED";
    FD1P3DX mem_9___i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_541), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[9] [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_9___i8.GSR = "ENABLED";
    FD1P3DX mem_9___i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_541), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[9] [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_9___i9.GSR = "ENABLED";
    FD1P3DX mem_9___i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_541), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[9] [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_9___i10.GSR = "ENABLED";
    FD1P3DX mem_9___i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_541), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[9] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_9___i11.GSR = "ENABLED";
    FD1P3DX mem_9___i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_541), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[9] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_9___i12.GSR = "ENABLED";
    FD1P3DX mem_9___i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_541), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[9] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_9___i13.GSR = "ENABLED";
    FD1P3DX mem_9___i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_541), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[9] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_9___i14.GSR = "ENABLED";
    FD1P3DX mem_9___i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_541), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[9] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_9___i15.GSR = "ENABLED";
    FD1P3BX mem_8___i2 (.D(din_reg[0]), .SP(REF_CLK_c_enable_556), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.smpl_width [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_8___i2.GSR = "ENABLED";
    FD1P3DX mem_8___i3 (.D(din_reg[1]), .SP(REF_CLK_c_enable_556), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[8] [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_8___i3.GSR = "ENABLED";
    FD1P3DX mem_8___i4 (.D(din_reg[2]), .SP(REF_CLK_c_enable_556), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[8] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_8___i4.GSR = "ENABLED";
    FD1P3DX mem_8___i5 (.D(din_reg[3]), .SP(REF_CLK_c_enable_556), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[8] [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_8___i5.GSR = "ENABLED";
    FD1P3DX mem_8___i6 (.D(din_reg[4]), .SP(REF_CLK_c_enable_556), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\inst2_from_fpgacfg.mode )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_8___i6.GSR = "ENABLED";
    FD1P3DX mem_8___i7 (.D(din_reg[5]), .SP(REF_CLK_c_enable_556), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\inst2_from_fpgacfg.ddr_en )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_8___i7.GSR = "ENABLED";
    FD1P3DX mem_8___i8 (.D(din_reg[6]), .SP(REF_CLK_c_enable_556), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\inst2_from_fpgacfg.trxiq_pulse )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_8___i8.GSR = "ENABLED";
    FD1P3BX mem_8___i9 (.D(din_reg[7]), .SP(REF_CLK_c_enable_556), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\inst2_from_fpgacfg.mimo_int_en )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_8___i9.GSR = "ENABLED";
    FD1P3DX mem_8___i10 (.D(din_reg[8]), .SP(REF_CLK_c_enable_556), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\inst2_from_fpgacfg.synch_dis )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_8___i10.GSR = "ENABLED";
    FD1P3DX mem_8___i11 (.D(din_reg[9]), .SP(REF_CLK_c_enable_556), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\inst2_from_fpgacfg.synch_mode )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_8___i11.GSR = "ENABLED";
    FD1P3DX mem_8___i12 (.D(din_reg[10]), .SP(REF_CLK_c_enable_556), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[8] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_8___i12.GSR = "ENABLED";
    FD1P3DX mem_8___i13 (.D(din_reg[11]), .SP(REF_CLK_c_enable_556), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[8] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_8___i13.GSR = "ENABLED";
    FD1P3DX mem_8___i14 (.D(din_reg[12]), .SP(REF_CLK_c_enable_556), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[8] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_8___i14.GSR = "ENABLED";
    FD1P3DX mem_8___i15 (.D(din_reg[13]), .SP(REF_CLK_c_enable_556), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[8] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_8___i15.GSR = "ENABLED";
    FD1P3DX mem_8___i16 (.D(din_reg[14]), .SP(REF_CLK_c_enable_556), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[8] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_8___i16.GSR = "ENABLED";
    FD1P3BX mem_7__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_571), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.ch_en [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_7__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_7__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_571), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.ch_en [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_7__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_7__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_571), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.ch_en [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_7__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_7__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_571), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.ch_en [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_7__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_7__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_571), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.ch_en [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_7__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_7__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_571), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.ch_en [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_7__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_7__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_571), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.ch_en [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_7__i0_i7.GSR = "ENABLED";
    FD1P3DX mem_7__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_571), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.ch_en [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_7__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_7__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_571), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.ch_en [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_7__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_7__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_571), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.ch_en [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_7__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_7__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_571), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.ch_en [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_7__i0_i11.GSR = "ENABLED";
    FD1P3DX mem_7__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_571), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.ch_en [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_7__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_7__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_571), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.ch_en [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_7__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_7__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_571), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.ch_en [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_7__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_7__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_571), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.ch_en [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_7__i0_i15.GSR = "ENABLED";
    FD1P3DX mem_6___i2 (.D(din_reg[0]), .SP(REF_CLK_c_enable_586), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.clk_ind [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_6___i2.GSR = "ENABLED";
    FD1P3DX mem_6___i3 (.D(din_reg[1]), .SP(REF_CLK_c_enable_586), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.clk_ind [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_6___i3.GSR = "ENABLED";
    FD1P3DX mem_6___i4 (.D(din_reg[2]), .SP(REF_CLK_c_enable_586), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.clk_ind [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_6___i4.GSR = "ENABLED";
    FD1P3DX mem_6___i5 (.D(din_reg[3]), .SP(REF_CLK_c_enable_586), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.clk_ind [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_6___i5.GSR = "ENABLED";
    FD1P3DX mem_6___i6 (.D(din_reg[4]), .SP(REF_CLK_c_enable_586), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.cnt_ind [0])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_6___i6.GSR = "ENABLED";
    FD1P3DX mem_6___i7 (.D(din_reg[5]), .SP(REF_CLK_c_enable_586), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.cnt_ind [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_6___i7.GSR = "ENABLED";
    FD1P3DX mem_6___i8 (.D(din_reg[6]), .SP(REF_CLK_c_enable_586), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.cnt_ind [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_6___i8.GSR = "ENABLED";
    FD1P3DX mem_6___i9 (.D(din_reg[7]), .SP(REF_CLK_c_enable_586), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.cnt_ind [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_6___i9.GSR = "ENABLED";
    FD1P3DX mem_6___i10 (.D(din_reg[8]), .SP(REF_CLK_c_enable_586), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.cnt_ind [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_6___i10.GSR = "ENABLED";
    FD1P3DX mem_6___i11 (.D(din_reg[9]), .SP(REF_CLK_c_enable_586), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\inst2_from_fpgacfg.load_phase_reg )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_6___i11.GSR = "ENABLED";
    FD1P3DX mem_6___i12 (.D(din_reg[10]), .SP(REF_CLK_c_enable_586), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[6] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_6___i12.GSR = "ENABLED";
    FD1P3DX mem_6___i13 (.D(din_reg[11]), .SP(REF_CLK_c_enable_586), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[6] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_6___i13.GSR = "ENABLED";
    FD1P3DX mem_6___i14 (.D(din_reg[12]), .SP(REF_CLK_c_enable_586), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[6] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_6___i14.GSR = "ENABLED";
    FD1P3DX mem_6___i15 (.D(din_reg[13]), .SP(REF_CLK_c_enable_586), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[6] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_6___i15.GSR = "ENABLED";
    FD1P3DX mem_6___i16 (.D(din_reg[14]), .SP(REF_CLK_c_enable_586), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[6] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_6___i16.GSR = "ENABLED";
    FD1P3DX mem_5__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_601), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.drct_clk_en [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_5__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_5__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_601), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.drct_clk_en [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_5__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_5__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_601), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.drct_clk_en [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_5__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_5__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_601), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.drct_clk_en [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_5__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_5__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_601), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.drct_clk_en [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_5__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_5__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_601), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.drct_clk_en [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_5__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_5__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_601), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.drct_clk_en [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_5__i0_i7.GSR = "ENABLED";
    FD1P3DX mem_5__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_601), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.drct_clk_en [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_5__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_5__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_601), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.drct_clk_en [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_5__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_5__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_601), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.drct_clk_en [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_5__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_5__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_601), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.drct_clk_en [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_5__i0_i11.GSR = "ENABLED";
    FD1P3DX mem_5__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_601), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.drct_clk_en [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_5__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_5__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_601), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.drct_clk_en [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_5__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_5__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_601), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.drct_clk_en [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_5__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_5__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_601), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.drct_clk_en [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_5__i0_i15.GSR = "ENABLED";
    FD1P3DX mem_4__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_616), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.phase_reg_sel [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_4__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_4__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_616), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.phase_reg_sel [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_4__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_4__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_616), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.phase_reg_sel [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_4__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_4__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_616), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.phase_reg_sel [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_4__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_4__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_616), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.phase_reg_sel [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_4__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_4__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_616), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.phase_reg_sel [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_4__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_4__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_616), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.phase_reg_sel [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_4__i0_i7.GSR = "ENABLED";
    FD1P3DX mem_4__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_616), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.phase_reg_sel [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_4__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_4__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_616), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.phase_reg_sel [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_4__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_4__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_616), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.phase_reg_sel [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_4__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_4__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_616), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.phase_reg_sel [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_4__i0_i11.GSR = "ENABLED";
    FD1P3DX mem_4__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_616), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.phase_reg_sel [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_4__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_4__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_616), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.phase_reg_sel [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_4__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_4__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_616), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.phase_reg_sel [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_4__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_4__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_616), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\from_fpgacfg.phase_reg_sel [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_4__i0_i15.GSR = "ENABLED";
    FD1P3DX mem_3__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_631), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[3] [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_3__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_3__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_631), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[3] [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_3__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_3__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_631), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[3] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_3__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_3__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_631), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[3] [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_3__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_3__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_631), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[3] [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_3__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_3__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_631), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[3] [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_3__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_3__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_631), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[3] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_3__i0_i7.GSR = "ENABLED";
    FD1P3DX mem_3__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_631), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[3] [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_3__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_3__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_631), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[3] [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_3__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_3__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_631), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[3] [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_3__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_3__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_631), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[3] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_3__i0_i11.GSR = "ENABLED";
    FD1P3DX mem_3__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_631), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[3] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_3__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_3__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_631), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[3] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_3__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_3__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_631), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[3] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_3__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_3__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_631), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[3] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_3__i0_i15.GSR = "ENABLED";
    FD1P3DX mem_2__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_646), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[2] [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_2__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_2__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_646), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[2] [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_2__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_2__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_646), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[2] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_2__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_2__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_646), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[2] [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_2__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_2__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_646), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[2] [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_2__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_2__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_646), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[2] [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_2__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_2__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_646), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[2] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_2__i0_i7.GSR = "ENABLED";
    FD1P3DX mem_2__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_646), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[2] [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_2__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_2__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_646), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[2] [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_2__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_2__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_646), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[2] [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_2__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_2__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_646), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[2] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_2__i0_i11.GSR = "ENABLED";
    FD1P3DX mem_2__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_646), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[2] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_2__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_2__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_646), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[2] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_2__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_2__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_646), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[2] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_2__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_2__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_646), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[2] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_2__i0_i15.GSR = "ENABLED";
    FD1P3DX mem_1__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_661), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[1] [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_1__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_1__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_661), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[1] [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_1__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_1__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_661), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[1] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_1__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_1__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_661), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[1] [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_1__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_1__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_661), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[1] [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_1__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_1__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_661), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[1] [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_1__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_1__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_661), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[1] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_1__i0_i7.GSR = "ENABLED";
    FD1P3DX mem_1__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_661), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[1] [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_1__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_1__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_661), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[1] [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_1__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_1__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_661), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[1] [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_1__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_1__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_661), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[1] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_1__i0_i11.GSR = "ENABLED";
    FD1P3DX mem_1__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_661), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[1] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_1__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_1__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_661), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[1] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_1__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_1__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_661), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[1] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_1__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_1__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_661), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[1] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_1__i0_i15.GSR = "ENABLED";
    FD1P3DX mem_0__i0_i1 (.D(din_reg[0]), .SP(REF_CLK_c_enable_676), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[0] [1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_0__i0_i1.GSR = "ENABLED";
    FD1P3DX mem_0__i0_i2 (.D(din_reg[1]), .SP(REF_CLK_c_enable_676), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[0] [2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_0__i0_i2.GSR = "ENABLED";
    FD1P3DX mem_0__i0_i3 (.D(din_reg[2]), .SP(REF_CLK_c_enable_676), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[0] [3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_0__i0_i3.GSR = "ENABLED";
    FD1P3DX mem_0__i0_i4 (.D(din_reg[3]), .SP(REF_CLK_c_enable_676), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[0] [4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_0__i0_i4.GSR = "ENABLED";
    FD1P3DX mem_0__i0_i5 (.D(din_reg[4]), .SP(REF_CLK_c_enable_676), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[0] [5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_0__i0_i5.GSR = "ENABLED";
    FD1P3DX mem_0__i0_i6 (.D(din_reg[5]), .SP(REF_CLK_c_enable_676), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[0] [6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_0__i0_i6.GSR = "ENABLED";
    FD1P3DX mem_0__i0_i7 (.D(din_reg[6]), .SP(REF_CLK_c_enable_676), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[0] [7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_0__i0_i7.GSR = "ENABLED";
    FD1P3DX mem_0__i0_i8 (.D(din_reg[7]), .SP(REF_CLK_c_enable_676), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[0] [8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_0__i0_i8.GSR = "ENABLED";
    FD1P3DX mem_0__i0_i9 (.D(din_reg[8]), .SP(REF_CLK_c_enable_676), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[0] [9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_0__i0_i9.GSR = "ENABLED";
    FD1P3DX mem_0__i0_i10 (.D(din_reg[9]), .SP(REF_CLK_c_enable_676), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[0] [10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_0__i0_i10.GSR = "ENABLED";
    FD1P3DX mem_0__i0_i11 (.D(din_reg[10]), .SP(REF_CLK_c_enable_676), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[0] [11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_0__i0_i11.GSR = "ENABLED";
    FD1P3DX mem_0__i0_i12 (.D(din_reg[11]), .SP(REF_CLK_c_enable_676), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[0] [12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_0__i0_i12.GSR = "ENABLED";
    FD1P3DX mem_0__i0_i13 (.D(din_reg[12]), .SP(REF_CLK_c_enable_676), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[0] [13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_0__i0_i13.GSR = "ENABLED";
    FD1P3DX mem_0__i0_i14 (.D(din_reg[13]), .SP(REF_CLK_c_enable_676), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[0] [14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_0__i0_i14.GSR = "ENABLED";
    FD1P3DX mem_0__i0_i15 (.D(din_reg[14]), .SP(REF_CLK_c_enable_676), .CK(REF_CLK_c), 
            .CD(n41434), .Q(\mem[0] [15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_0__i0_i15.GSR = "ENABLED";
    L6MUX21 i32153 (.D0(n37323), .D1(n37324), .SD(inst_reg[2]), .Z(n37325));
    L6MUX21 i32160 (.D0(n37330), .D1(n37331), .SD(inst_reg[2]), .Z(n37332));
    L6MUX21 i32167 (.D0(n37337), .D1(n37338), .SD(inst_reg[2]), .Z(n37339));
    L6MUX21 i32174 (.D0(n37344), .D1(n37345), .SD(inst_reg[2]), .Z(n37346));
    LUT4 i32026_3_lut_4_lut_then_4_lut (.A(inst_reg[1]), .B(inst_reg[2]), 
         .C(\mem[24] [3]), .D(\mem[26] [3]), .Z(n41454)) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam i32026_3_lut_4_lut_then_4_lut.init = 16'hc480;
    L6MUX21 i32181 (.D0(n37351), .D1(n37352), .SD(inst_reg[2]), .Z(n37353));
    LUT4 i31136_3_lut (.A(\mem[25] [13]), .B(\mem[24] [13]), .C(inst_reg[0]), 
         .Z(n36308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31136_3_lut.init = 16'hcaca;
    L6MUX21 i32188 (.D0(n37358), .D1(n37359), .SD(inst_reg[2]), .Z(n37360));
    L6MUX21 i32195 (.D0(n37365), .D1(n37366), .SD(inst_reg[2]), .Z(n37367));
    L6MUX21 i32202 (.D0(n37372), .D1(n37373), .SD(inst_reg[2]), .Z(n37374));
    L6MUX21 i32209 (.D0(n37379), .D1(n37380), .SD(inst_reg[2]), .Z(n37381));
    L6MUX21 i32216 (.D0(n37386), .D1(n37387), .SD(inst_reg[2]), .Z(n37388));
    L6MUX21 i32223 (.D0(n37393), .D1(n37394), .SD(inst_reg[2]), .Z(n37395));
    L6MUX21 i32230 (.D0(n37400), .D1(n37401), .SD(inst_reg[2]), .Z(n37402));
    L6MUX21 i32237 (.D0(n37407), .D1(n37408), .SD(inst_reg[2]), .Z(n37409));
    L6MUX21 i32244 (.D0(n37414), .D1(n37415), .SD(inst_reg[2]), .Z(n37416));
    L6MUX21 i32251 (.D0(n37421), .D1(n37422), .SD(inst_reg[2]), .Z(n37423));
    LUT4 i31135_3_lut (.A(\mem[27] [13]), .B(\mem[26] [13]), .C(inst_reg[0]), 
         .Z(n36307)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31135_3_lut.init = 16'hcaca;
    L6MUX21 i32258 (.D0(n37428), .D1(n37429), .SD(inst_reg[2]), .Z(n37430));
    L6MUX21 i32265 (.D0(n37435), .D1(n37436), .SD(inst_reg[2]), .Z(n37437));
    L6MUX21 i32272 (.D0(n37442), .D1(n37443), .SD(inst_reg[2]), .Z(n37444));
    L6MUX21 i32279 (.D0(n37449), .D1(n37450), .SD(inst_reg[2]), .Z(n37451));
    L6MUX21 i32286 (.D0(n37456), .D1(n37457), .SD(inst_reg[2]), .Z(n37458));
    LUT4 i31133_3_lut (.A(\mem[25] [14]), .B(\mem[24] [14]), .C(inst_reg[0]), 
         .Z(n36305)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31133_3_lut.init = 16'hcaca;
    L6MUX21 i32293 (.D0(n37463), .D1(n37464), .SD(inst_reg[2]), .Z(n37465));
    L6MUX21 i32300 (.D0(n37470), .D1(n37471), .SD(inst_reg[2]), .Z(n37472));
    PFUMX i32309 (.BLUT(n37473), .ALUT(n37474), .C0(inst_reg[2]), .Z(n37481));
    LUT4 i31132_3_lut (.A(\mem[27] [14]), .B(\mem[26] [14]), .C(inst_reg[0]), 
         .Z(n36304)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31132_3_lut.init = 16'hcaca;
    LUT4 i31121_3_lut (.A(\mem[25] [15]), .B(\mem[24] [15]), .C(inst_reg[0]), 
         .Z(n36293)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31121_3_lut.init = 16'hcaca;
    LUT4 i31120_3_lut (.A(\mem[27] [15]), .B(\mem[26] [15]), .C(inst_reg[0]), 
         .Z(n36292)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31120_3_lut.init = 16'hcaca;
    L6MUX21 i32310 (.D0(n37475), .D1(n37476), .SD(inst_reg[2]), .Z(n37482));
    L6MUX21 i32311 (.D0(n37477), .D1(n37478), .SD(inst_reg[2]), .Z(n37483));
    L6MUX21 i32312 (.D0(n37479), .D1(n37480), .SD(inst_reg[2]), .Z(n37484));
    L6MUX21 i32317 (.D0(n36168), .D1(n36165), .SD(inst_reg[2]), .Z(n37489));
    L6MUX21 i32318 (.D0(n36162), .D1(n36159), .SD(inst_reg[2]), .Z(n37490));
    L6MUX21 i32319 (.D0(n36156), .D1(n36153), .SD(inst_reg[2]), .Z(n37491));
    LUT4 i30875_3_lut (.A(\mem[1] [1]), .B(\mem[0] [1]), .C(inst_reg[0]), 
         .Z(n36047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30875_3_lut.init = 16'hcaca;
    LUT4 i30874_3_lut (.A(\mem[3] [1]), .B(\mem[2] [1]), .C(inst_reg[0]), 
         .Z(n36046)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30874_3_lut.init = 16'hcaca;
    LUT4 i30872_3_lut (.A(\from_fpgacfg.drct_clk_en [1]), .B(\from_fpgacfg.phase_reg_sel [1]), 
         .C(inst_reg[0]), .Z(n36044)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30872_3_lut.init = 16'hcaca;
    LUT4 i32322_3_lut (.A(n37492), .B(n37493), .C(inst_reg[4]), .Z(dout_reg_15__N_5274[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32322_3_lut.init = 16'hcaca;
    LUT4 i30871_3_lut (.A(\from_fpgacfg.ch_en [1]), .B(\from_fpgacfg.clk_ind [1]), 
         .C(inst_reg[0]), .Z(n36043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30871_3_lut.init = 16'hcaca;
    LUT4 i30869_3_lut (.A(\inst2_from_fpgacfg.txpct_loss_clr ), .B(\from_fpgacfg.smpl_width [1]), 
         .C(inst_reg[0]), .Z(n36041)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30869_3_lut.init = 16'hcaca;
    LUT4 i30868_3_lut (.A(\mem[11] [1]), .B(\inst2_from_fpgacfg.tx_en ), 
         .C(inst_reg[0]), .Z(n36040)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30868_3_lut.init = 16'hcaca;
    LUT4 i30866_3_lut (.A(\inst2_from_fpgacfg.wfm_play ), .B(\from_fpgacfg.wfm_ch_en [1]), 
         .C(inst_reg[0]), .Z(n36038)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30866_3_lut.init = 16'hcaca;
    LUT4 i30865_3_lut (.A(\from_fpgacfg.sync_size [1]), .B(\mem[14] [1]), 
         .C(inst_reg[0]), .Z(n36037)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30865_3_lut.init = 16'hcaca;
    LUT4 i30863_3_lut (.A(\from_fpgacfg.txant_post [1]), .B(\from_fpgacfg.txant_pre [1]), 
         .C(inst_reg[0]), .Z(n36035)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30863_3_lut.init = 16'hcaca;
    LUT4 i30862_3_lut (.A(\inst2_from_fpgacfg.LMS1_RESET ), .B(\mem[18] [1]), 
         .C(inst_reg[0]), .Z(n36034)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30862_3_lut.init = 16'hcaca;
    LUT4 i30860_3_lut (.A(\mem[21] [1]), .B(\mem[20] [1]), .C(inst_reg[0]), 
         .Z(n36032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30860_3_lut.init = 16'hcaca;
    LUT4 i30859_3_lut (.A(\from_fpgacfg.GPIO [1]), .B(\mem[22] [1]), .C(inst_reg[0]), 
         .Z(n36031)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30859_3_lut.init = 16'hcaca;
    LUT4 i32320_3_lut (.A(n37488), .B(n37489), .C(inst_reg[3]), .Z(n37492)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32320_3_lut.init = 16'hcaca;
    LUT4 i32316_4_lut (.A(n41431), .B(n36174), .C(inst_reg[2]), .D(hw_ver_int[2]), 
         .Z(n37488)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;
    defparam i32316_4_lut.init = 16'hcfc5;
    LUT4 i30851_3_lut (.A(\mem[1] [3]), .B(\mem[0] [3]), .C(inst_reg[0]), 
         .Z(n36023)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30851_3_lut.init = 16'hcaca;
    LUT4 i30850_3_lut (.A(\mem[3] [3]), .B(\mem[2] [3]), .C(inst_reg[0]), 
         .Z(n36022)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30850_3_lut.init = 16'hcaca;
    LUT4 i32025_3_lut (.A(n37195), .B(n37196), .C(inst_reg[4]), .Z(dout_reg_15__N_5274[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32025_3_lut.init = 16'hcaca;
    LUT4 i32023_3_lut (.A(n37191), .B(n37192), .C(inst_reg[3]), .Z(n37195)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32023_3_lut.init = 16'hcaca;
    LUT4 i32019_4_lut (.A(n20513), .B(n35982), .C(inst_reg[2]), .D(inst_reg[0]), 
         .Z(n37191)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;
    defparam i32019_4_lut.init = 16'hcacf;
    LUT4 i15247_2_lut (.A(inst_reg[1]), .B(hw_ver_int[2]), .Z(n20513)) /* synthesis lut_function=(A (B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam i15247_2_lut.init = 16'h8888;
    LUT4 i32032_3_lut (.A(n37202), .B(n37203), .C(inst_reg[4]), .Z(dout_reg_15__N_5274[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32032_3_lut.init = 16'hcaca;
    LUT4 i32030_3_lut (.A(n41455), .B(n37199), .C(inst_reg[3]), .Z(n37202)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32030_3_lut.init = 16'hcaca;
    LUT4 i32315_3_lut (.A(n37485), .B(n37486), .C(inst_reg[4]), .Z(dout_reg_15__N_5274[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32315_3_lut.init = 16'hcaca;
    LUT4 i30848_3_lut (.A(\from_fpgacfg.drct_clk_en [3]), .B(\from_fpgacfg.phase_reg_sel [3]), 
         .C(inst_reg[0]), .Z(n36020)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30848_3_lut.init = 16'hcaca;
    LUT4 i30847_3_lut (.A(\from_fpgacfg.ch_en [3]), .B(\from_fpgacfg.clk_ind [3]), 
         .C(inst_reg[0]), .Z(n36019)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30847_3_lut.init = 16'hcaca;
    LUT4 i32313_3_lut (.A(n37481), .B(n37482), .C(inst_reg[3]), .Z(n37485)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32313_3_lut.init = 16'hcaca;
    LUT4 i30845_3_lut (.A(\mem[9] [3]), .B(\mem[8] [3]), .C(inst_reg[0]), 
         .Z(n36017)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30845_3_lut.init = 16'hcaca;
    LUT4 i32039_3_lut (.A(n37209), .B(n37210), .C(inst_reg[4]), .Z(dout_reg_15__N_5274[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32039_3_lut.init = 16'hcaca;
    LUT4 i32037_3_lut (.A(n41458), .B(n37206), .C(inst_reg[3]), .Z(n37209)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32037_3_lut.init = 16'hcaca;
    LUT4 i30844_3_lut (.A(\mem[11] [3]), .B(\mem[10] [3]), .C(inst_reg[0]), 
         .Z(n36016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30844_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n1800[31]), .B(n41191), .C(n11789), 
         .D(n41446), .Z(REF_CLK_c_enable_367)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1010 (.A(n1800[31]), .B(n41191), .C(n30140), 
         .D(n41446), .Z(REF_CLK_c_enable_304)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1010.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1011 (.A(n1800[31]), .B(n41191), .C(n31780), 
         .D(n41446), .Z(REF_CLK_c_enable_242)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1011.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1012 (.A(n1800[31]), .B(n41191), .C(n31786), 
         .D(n41446), .Z(REF_CLK_c_enable_526)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1012.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1013 (.A(n1800[31]), .B(n41191), .C(n30139), 
         .D(n41446), .Z(REF_CLK_c_enable_586)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1013.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1014 (.A(n1800[31]), .B(n41191), .C(n11264), 
         .D(n41446), .Z(REF_CLK_c_enable_1608)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1014.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1015 (.A(n1800[31]), .B(n41191), .C(n11789), 
         .D(n41431), .Z(REF_CLK_c_enable_382)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1015.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1016 (.A(n1800[31]), .B(n41191), .C(n30140), 
         .D(n41431), .Z(REF_CLK_c_enable_322)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1016.init = 16'h0800;
    LUT4 mux_16_Mux_2_i24_3_lut (.A(\from_fpgacfg.drct_clk_en [2]), .B(\from_fpgacfg.phase_reg_sel [2]), 
         .C(inst_reg[0]), .Z(n24)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam mux_16_Mux_2_i24_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1017 (.A(n1800[31]), .B(n41191), .C(n31780), 
         .D(n41431), .Z(REF_CLK_c_enable_258)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1017.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1018 (.A(n1800[31]), .B(n41191), .C(n31786), 
         .D(n41431), .Z(REF_CLK_c_enable_511)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1018.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1019 (.A(n1800[31]), .B(n41191), .C(n30139), 
         .D(n41431), .Z(REF_CLK_c_enable_571)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1019.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1020 (.A(n1800[31]), .B(n41191), .C(n11264), 
         .D(n41431), .Z(REF_CLK_c_enable_202)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1020.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1021 (.A(n1800[31]), .B(n41191), .C(n11264), 
         .D(n41384), .Z(REF_CLK_c_enable_384)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1021.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1022 (.A(n1800[31]), .B(n41191), .C(n11789), 
         .D(n41384), .Z(REF_CLK_c_enable_337)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1022.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1023 (.A(n1800[31]), .B(n41191), .C(n30140), 
         .D(n41384), .Z(REF_CLK_c_enable_273)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1023.init = 16'h0008;
    PFUMX i30789 (.BLUT(n35959), .ALUT(n35960), .C0(inst_reg[1]), .Z(n35961));
    LUT4 i1_2_lut_3_lut_4_lut_adj_1024 (.A(n1800[31]), .B(n41191), .C(n31780), 
         .D(n41384), .Z(REF_CLK_c_enable_211)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1024.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1025 (.A(n1800[31]), .B(n41191), .C(n31786), 
         .D(n41384), .Z(REF_CLK_c_enable_556)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1025.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1026 (.A(n1800[31]), .B(n41191), .C(n30139), 
         .D(n41384), .Z(REF_CLK_c_enable_616)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1026.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1027 (.A(n1800[31]), .B(n41191), .C(n11264), 
         .D(n41447), .Z(REF_CLK_c_enable_387)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1027.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1028 (.A(n1800[31]), .B(n41191), .C(n11789), 
         .D(n41447), .Z(REF_CLK_c_enable_352)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1028.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1029 (.A(n1800[31]), .B(n41191), .C(n30140), 
         .D(n41447), .Z(REF_CLK_c_enable_289)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1029.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1030 (.A(n1800[31]), .B(n41191), .C(n31780), 
         .D(n41447), .Z(REF_CLK_c_enable_226)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1030.init = 16'h0008;
    PFUMX i30792 (.BLUT(n35962), .ALUT(n35963), .C0(inst_reg[1]), .Z(n35964));
    LUT4 mux_16_Mux_2_i23_3_lut (.A(\from_fpgacfg.ch_en [2]), .B(\from_fpgacfg.clk_ind [2]), 
         .C(inst_reg[0]), .Z(n23)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam mux_16_Mux_2_i23_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1031 (.A(n1800[31]), .B(n41191), .C(n31786), 
         .D(n41447), .Z(REF_CLK_c_enable_541)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1031.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1032 (.A(n1800[31]), .B(n41191), .C(n30139), 
         .D(n41447), .Z(REF_CLK_c_enable_601)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1032.init = 16'h0008;
    LUT4 i1_2_lut_rep_769_3_lut (.A(n1800[31]), .B(n41191), .C(inst_reg[4]), 
         .Z(n41174)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_769_3_lut.init = 16'h0808;
    LUT4 i31102_4_lut (.A(n36294), .B(n37248), .C(inst_reg[3]), .D(inst_reg[2]), 
         .Z(n36274)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i31102_4_lut.init = 16'hcac0;
    LUT4 i31129_4_lut (.A(n36306), .B(n37269), .C(inst_reg[3]), .D(inst_reg[2]), 
         .Z(n36301)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i31129_4_lut.init = 16'hcac0;
    LUT4 i31138_4_lut (.A(n36309), .B(n37290), .C(inst_reg[3]), .D(inst_reg[2]), 
         .Z(n36310)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i31138_4_lut.init = 16'hcac0;
    LUT4 i30784_4_lut (.A(n36315), .B(n37311), .C(inst_reg[3]), .D(inst_reg[2]), 
         .Z(n35956)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i30784_4_lut.init = 16'hcac0;
    LUT4 i30838_4_lut (.A(n35961), .B(n37332), .C(inst_reg[3]), .D(inst_reg[2]), 
         .Z(n36010)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i30838_4_lut.init = 16'hcac0;
    LUT4 i30853_4_lut (.A(n35964), .B(n37353), .C(inst_reg[3]), .D(inst_reg[2]), 
         .Z(n36025)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i30853_4_lut.init = 16'hcac0;
    LUT4 i31114_4_lut (.A(n35967), .B(n37374), .C(inst_reg[3]), .D(inst_reg[2]), 
         .Z(n36286)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i31114_4_lut.init = 16'hcac0;
    PFUMX i30795 (.BLUT(n35965), .ALUT(n35966), .C0(inst_reg[1]), .Z(n35967));
    LUT4 i31117_4_lut (.A(n35970), .B(n37395), .C(inst_reg[3]), .D(inst_reg[2]), 
         .Z(n36289)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i31117_4_lut.init = 16'hcac0;
    LUT4 i31123_4_lut (.A(n35973), .B(n37416), .C(inst_reg[3]), .D(inst_reg[2]), 
         .Z(n36295)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i31123_4_lut.init = 16'hcac0;
    LUT4 i31126_4_lut (.A(n35976), .B(n37437), .C(inst_reg[3]), .D(inst_reg[2]), 
         .Z(n36298)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i31126_4_lut.init = 16'hcac0;
    LUT4 i30877_4_lut (.A(n35979), .B(n37458), .C(inst_reg[3]), .D(inst_reg[2]), 
         .Z(n36049)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i30877_4_lut.init = 16'hcac0;
    PFUMX i30798 (.BLUT(n35968), .ALUT(n35969), .C0(inst_reg[1]), .Z(n35970));
    PFUMX i30801 (.BLUT(n35971), .ALUT(n35972), .C0(inst_reg[1]), .Z(n35973));
    PFUMX i30804 (.BLUT(n35974), .ALUT(n35975), .C0(inst_reg[1]), .Z(n35976));
    PFUMX i30807 (.BLUT(n35977), .ALUT(n35978), .C0(inst_reg[1]), .Z(n35979));
    FD1P3DX inst_reg_i0_i1 (.D(inst_reg[0]), .SP(REF_CLK_c_enable_1424), 
            .CK(REF_CLK_c), .CD(n41434), .Q(inst_reg[1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(115[7] 124[14])
    defparam inst_reg_i0_i1.GSR = "ENABLED";
    FD1P3DX inst_reg_i0_i2 (.D(inst_reg[1]), .SP(REF_CLK_c_enable_1424), 
            .CK(REF_CLK_c), .CD(n41434), .Q(inst_reg[2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(115[7] 124[14])
    defparam inst_reg_i0_i2.GSR = "ENABLED";
    FD1P3DX inst_reg_i0_i3 (.D(inst_reg[2]), .SP(REF_CLK_c_enable_1424), 
            .CK(REF_CLK_c), .CD(n41434), .Q(inst_reg[3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(115[7] 124[14])
    defparam inst_reg_i0_i3.GSR = "ENABLED";
    FD1P3DX inst_reg_i0_i4 (.D(inst_reg[3]), .SP(REF_CLK_c_enable_1424), 
            .CK(REF_CLK_c), .CD(n41434), .Q(inst_reg[4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(115[7] 124[14])
    defparam inst_reg_i0_i4.GSR = "ENABLED";
    FD1P3DX inst_reg_i0_i5 (.D(inst_reg[4]), .SP(REF_CLK_c_enable_1424), 
            .CK(REF_CLK_c), .CD(n41434), .Q(inst_reg[5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(115[7] 124[14])
    defparam inst_reg_i0_i5.GSR = "ENABLED";
    FD1P3DX inst_reg_i0_i6 (.D(inst_reg[5]), .SP(REF_CLK_c_enable_1424), 
            .CK(REF_CLK_c), .CD(n41434), .Q(inst_reg[6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(115[7] 124[14])
    defparam inst_reg_i0_i6.GSR = "ENABLED";
    FD1P3DX inst_reg_i0_i7 (.D(inst_reg[6]), .SP(REF_CLK_c_enable_1424), 
            .CK(REF_CLK_c), .CD(n41434), .Q(inst_reg[7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(115[7] 124[14])
    defparam inst_reg_i0_i7.GSR = "ENABLED";
    FD1P3DX inst_reg_i0_i8 (.D(inst_reg[7]), .SP(REF_CLK_c_enable_1424), 
            .CK(REF_CLK_c), .CD(n41434), .Q(inst_reg[8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(115[7] 124[14])
    defparam inst_reg_i0_i8.GSR = "ENABLED";
    FD1P3DX inst_reg_i0_i9 (.D(inst_reg[8]), .SP(REF_CLK_c_enable_1424), 
            .CK(REF_CLK_c), .CD(n41434), .Q(inst_reg[9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(115[7] 124[14])
    defparam inst_reg_i0_i9.GSR = "ENABLED";
    FD1P3DX inst_reg_i0_i10 (.D(inst_reg[9]), .SP(REF_CLK_c_enable_1424), 
            .CK(REF_CLK_c), .CD(n41434), .Q(inst_reg[10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(115[7] 124[14])
    defparam inst_reg_i0_i10.GSR = "ENABLED";
    FD1P3DX inst_reg_i0_i11 (.D(inst_reg[10]), .SP(REF_CLK_c_enable_1424), 
            .CK(REF_CLK_c), .CD(n41434), .Q(inst_reg[11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(115[7] 124[14])
    defparam inst_reg_i0_i11.GSR = "ENABLED";
    FD1P3DX inst_reg_i0_i12 (.D(inst_reg[11]), .SP(REF_CLK_c_enable_1424), 
            .CK(REF_CLK_c), .CD(n41434), .Q(inst_reg[12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(115[7] 124[14])
    defparam inst_reg_i0_i12.GSR = "ENABLED";
    FD1P3DX inst_reg_i0_i13 (.D(inst_reg[12]), .SP(REF_CLK_c_enable_1424), 
            .CK(REF_CLK_c), .CD(n41434), .Q(inst_reg[13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(115[7] 124[14])
    defparam inst_reg_i0_i13.GSR = "ENABLED";
    FD1P3DX inst_reg_i0_i14 (.D(inst_reg[13]), .SP(REF_CLK_c_enable_1424), 
            .CK(REF_CLK_c), .CD(n41434), .Q(inst_reg[14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(115[7] 124[14])
    defparam inst_reg_i0_i14.GSR = "ENABLED";
    FD1P3DX inst_reg_i0_i15 (.D(inst_reg[14]), .SP(REF_CLK_c_enable_1424), 
            .CK(REF_CLK_c), .CD(n41434), .Q(\inst_reg[15] )) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(115[7] 124[14])
    defparam inst_reg_i0_i15.GSR = "ENABLED";
    LUT4 mux_16_Mux_2_i20_3_lut (.A(\mem[9] [2]), .B(\mem[8] [2]), .C(inst_reg[0]), 
         .Z(n20)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam mux_16_Mux_2_i20_3_lut.init = 16'hcaca;
    LUT4 mux_16_Mux_2_i19_3_lut (.A(\mem[11] [2]), .B(\mem[10] [2]), .C(inst_reg[0]), 
         .Z(n19)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam mux_16_Mux_2_i19_3_lut.init = 16'hcaca;
    LUT4 mux_16_Mux_2_i17_3_lut (.A(\inst2_from_fpgacfg.wfm_load ), .B(\from_fpgacfg.wfm_ch_en [2]), 
         .C(inst_reg[0]), .Z(n17)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam mux_16_Mux_2_i17_3_lut.init = 16'hcaca;
    PFUMX i30810 (.BLUT(n35980), .ALUT(n35981), .C0(inst_reg[1]), .Z(n35982));
    PFUMX i30813 (.BLUT(n35983), .ALUT(n35984), .C0(inst_reg[1]), .Z(n35985));
    LUT4 i30842_3_lut (.A(\mem[13] [3]), .B(\from_fpgacfg.wfm_ch_en [3]), 
         .C(inst_reg[0]), .Z(n36014)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30842_3_lut.init = 16'hcaca;
    PFUMX i30816 (.BLUT(n35986), .ALUT(n35987), .C0(inst_reg[1]), .Z(n35988));
    PFUMX i30819 (.BLUT(n35989), .ALUT(n35990), .C0(inst_reg[1]), .Z(n35991));
    PFUMX i30822 (.BLUT(n35992), .ALUT(n35993), .C0(inst_reg[1]), .Z(n35994));
    PFUMX i30825 (.BLUT(n35995), .ALUT(n35996), .C0(inst_reg[1]), .Z(n35997));
    PFUMX i30828 (.BLUT(n35998), .ALUT(n35999), .C0(inst_reg[1]), .Z(n36000));
    LUT4 i30841_3_lut (.A(\from_fpgacfg.sync_size [3]), .B(\mem[14] [3]), 
         .C(inst_reg[0]), .Z(n36013)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30841_3_lut.init = 16'hcaca;
    LUT4 i30836_3_lut (.A(\from_fpgacfg.txant_post [3]), .B(\from_fpgacfg.txant_pre [3]), 
         .C(inst_reg[0]), .Z(n36008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30836_3_lut.init = 16'hcaca;
    LUT4 mux_16_Mux_2_i16_3_lut (.A(\from_fpgacfg.sync_size [2]), .B(\mem[14] [2]), 
         .C(inst_reg[0]), .Z(n16)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam mux_16_Mux_2_i16_3_lut.init = 16'hcaca;
    LUT4 mux_16_Mux_2_i12_3_lut (.A(\from_fpgacfg.txant_post [2]), .B(\from_fpgacfg.txant_pre [2]), 
         .C(inst_reg[0]), .Z(n12)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam mux_16_Mux_2_i12_3_lut.init = 16'hcaca;
    PFUMX i30834 (.BLUT(n36004), .ALUT(n36005), .C0(inst_reg[1]), .Z(n36006));
    LUT4 i30835_3_lut (.A(\inst2_from_fpgacfg.LMS1_TXNRX1 ), .B(\mem[18] [3]), 
         .C(inst_reg[0]), .Z(n36007)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30835_3_lut.init = 16'hcaca;
    LUT4 i30833_3_lut (.A(\mem[21] [3]), .B(\mem[20] [3]), .C(inst_reg[0]), 
         .Z(n36005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30833_3_lut.init = 16'hcaca;
    LUT4 i30832_3_lut (.A(\from_fpgacfg.GPIO [3]), .B(\mem[22] [3]), .C(inst_reg[0]), 
         .Z(n36004)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30832_3_lut.init = 16'hcaca;
    PFUMX i30837 (.BLUT(n36007), .ALUT(n36008), .C0(inst_reg[1]), .Z(n36009));
    FD1P3DX din_reg__i2 (.D(din_reg[0]), .SP(REF_CLK_c_enable_1621), .CK(REF_CLK_c), 
            .CD(n41434), .Q(din_reg[1])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(133[7] 142[14])
    defparam din_reg__i2.GSR = "ENABLED";
    LUT4 mux_16_Mux_2_i11_3_lut (.A(\inst2_from_fpgacfg.LMS1_CORE_LDO_EN ), 
         .B(\mem[18] [2]), .C(inst_reg[0]), .Z(n11)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam mux_16_Mux_2_i11_3_lut.init = 16'hcaca;
    LUT4 mux_16_Mux_2_i9_3_lut (.A(\mem[21] [2]), .B(\mem[20] [2]), .C(inst_reg[0]), 
         .Z(n9)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam mux_16_Mux_2_i9_3_lut.init = 16'hcaca;
    LUT4 mux_16_Mux_2_i8_3_lut (.A(\from_fpgacfg.GPIO [2]), .B(\mem[22] [2]), 
         .C(inst_reg[0]), .Z(n8)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam mux_16_Mux_2_i8_3_lut.init = 16'hcaca;
    LUT4 mux_16_Mux_2_i5_3_lut (.A(\mem[25] [2]), .B(\mem[24] [2]), .C(inst_reg[0]), 
         .Z(n5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam mux_16_Mux_2_i5_3_lut.init = 16'hcaca;
    PFUMX i30843 (.BLUT(n36013), .ALUT(n36014), .C0(inst_reg[1]), .Z(n36015));
    FD1P3BX mem_30___i1 (.D(IO_MOSI_c), .SP(REF_CLK_c_enable_1608), .CK(REF_CLK_c), 
            .PD(n41434), .Q(\from_fpgacfg.sync_pulse_period [16])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(213[7] 262[14])
    defparam mem_30___i1.GSR = "ENABLED";
    LUT4 i30827_3_lut (.A(\mem[1] [4]), .B(\mem[0] [4]), .C(inst_reg[0]), 
         .Z(n35999)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30827_3_lut.init = 16'hcaca;
    LUT4 mux_16_Mux_2_i4_3_lut (.A(\mem[27] [2]), .B(\from_fpgacfg.FPGA_LED1_CTRL [2]), 
         .C(inst_reg[0]), .Z(n4)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam mux_16_Mux_2_i4_3_lut.init = 16'hcaca;
    LUT4 i32472_3_lut (.A(n4), .B(n5), .C(inst_reg[1]), .Z(n37474)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32472_3_lut.init = 16'hcaca;
    LUT4 i30826_3_lut (.A(\mem[3] [4]), .B(\mem[2] [4]), .C(inst_reg[0]), 
         .Z(n35998)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30826_3_lut.init = 16'hcaca;
    LUT4 i30824_3_lut (.A(\from_fpgacfg.drct_clk_en [4]), .B(\from_fpgacfg.phase_reg_sel [4]), 
         .C(inst_reg[0]), .Z(n35996)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30824_3_lut.init = 16'hcaca;
    LUT4 i30823_3_lut (.A(\from_fpgacfg.ch_en [4]), .B(\from_fpgacfg.clk_ind [4]), 
         .C(inst_reg[0]), .Z(n35995)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30823_3_lut.init = 16'hcaca;
    PFUMX i30846 (.BLUT(n36016), .ALUT(n36017), .C0(inst_reg[1]), .Z(n36018));
    LUT4 i30821_3_lut (.A(\mem[9] [4]), .B(\mem[8] [4]), .C(inst_reg[0]), 
         .Z(n35993)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30821_3_lut.init = 16'hcaca;
    LUT4 i30820_3_lut (.A(\mem[11] [4]), .B(\mem[10] [4]), .C(inst_reg[0]), 
         .Z(n35992)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30820_3_lut.init = 16'hcaca;
    LUT4 i30818_3_lut (.A(\mem[13] [4]), .B(\from_fpgacfg.wfm_ch_en [4]), 
         .C(inst_reg[0]), .Z(n35990)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30818_3_lut.init = 16'hcaca;
    LUT4 i30817_3_lut (.A(\from_fpgacfg.sync_size [4]), .B(\mem[14] [4]), 
         .C(inst_reg[0]), .Z(n35989)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30817_3_lut.init = 16'hcaca;
    LUT4 i30815_3_lut (.A(\from_fpgacfg.txant_post [4]), .B(\from_fpgacfg.txant_pre [4]), 
         .C(inst_reg[0]), .Z(n35987)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30815_3_lut.init = 16'hcaca;
    LUT4 i30814_3_lut (.A(\inst2_from_fpgacfg.LMS1_TXNRX2 ), .B(\mem[18] [4]), 
         .C(inst_reg[0]), .Z(n35986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30814_3_lut.init = 16'hcaca;
    LUT4 i30812_3_lut (.A(\mem[21] [4]), .B(\mem[20] [4]), .C(inst_reg[0]), 
         .Z(n35984)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30812_3_lut.init = 16'hcaca;
    LUT4 i30811_3_lut (.A(\from_fpgacfg.GPIO [4]), .B(\mem[22] [4]), .C(inst_reg[0]), 
         .Z(n35983)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30811_3_lut.init = 16'hcaca;
    LUT4 i30809_3_lut (.A(\mem[25] [4]), .B(\mem[24] [4]), .C(inst_reg[0]), 
         .Z(n35981)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30809_3_lut.init = 16'hcaca;
    LUT4 i30808_3_lut (.A(\mem[27] [4]), .B(\from_fpgacfg.FPGA_LED2_CTRL [0]), 
         .C(inst_reg[0]), .Z(n35980)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30808_3_lut.init = 16'hcaca;
    LUT4 i31001_3_lut (.A(\mem[25] [0]), .B(\mem[24] [0]), .C(inst_reg[0]), 
         .Z(n36173)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31001_3_lut.init = 16'hcaca;
    LUT4 i30806_3_lut (.A(\mem[25] [5]), .B(\mem[24] [5]), .C(inst_reg[0]), 
         .Z(n35978)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30806_3_lut.init = 16'hcaca;
    LUT4 i30805_3_lut (.A(\mem[27] [5]), .B(\from_fpgacfg.FPGA_LED2_CTRL [1]), 
         .C(inst_reg[0]), .Z(n35977)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30805_3_lut.init = 16'hcaca;
    LUT4 i30803_3_lut (.A(\mem[25] [6]), .B(\mem[24] [6]), .C(inst_reg[0]), 
         .Z(n35975)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30803_3_lut.init = 16'hcaca;
    LUT4 i31000_3_lut (.A(\mem[27] [0]), .B(\from_fpgacfg.FPGA_LED1_CTRL [0]), 
         .C(inst_reg[0]), .Z(n36172)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31000_3_lut.init = 16'hcaca;
    LUT4 i30802_3_lut (.A(\mem[27] [6]), .B(\from_fpgacfg.FPGA_LED2_CTRL [2]), 
         .C(inst_reg[0]), .Z(n35974)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30802_3_lut.init = 16'hcaca;
    LUT4 i30800_3_lut (.A(\mem[25] [7]), .B(\mem[24] [7]), .C(inst_reg[0]), 
         .Z(n35972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30800_3_lut.init = 16'hcaca;
    LUT4 i30799_3_lut (.A(\mem[27] [7]), .B(\mem[26] [7]), .C(inst_reg[0]), 
         .Z(n35971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30799_3_lut.init = 16'hcaca;
    LUT4 i30995_3_lut (.A(\mem[21] [0]), .B(\mem[20] [0]), .C(inst_reg[0]), 
         .Z(n36167)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30995_3_lut.init = 16'hcaca;
    LUT4 i30797_3_lut (.A(\mem[25] [8]), .B(\mem[24] [8]), .C(inst_reg[0]), 
         .Z(n35969)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30797_3_lut.init = 16'hcaca;
    LUT4 i30796_3_lut (.A(\mem[27] [8]), .B(\mem[26] [8]), .C(inst_reg[0]), 
         .Z(n35968)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30796_3_lut.init = 16'hcaca;
    LUT4 i30794_3_lut (.A(\mem[25] [9]), .B(\mem[24] [9]), .C(inst_reg[0]), 
         .Z(n35966)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30794_3_lut.init = 16'hcaca;
    LUT4 equal_240_i6_2_lut_rep_979 (.A(inst_reg[0]), .B(inst_reg[1]), .Z(n41384)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(253[20:62])
    defparam equal_240_i6_2_lut_rep_979.init = 16'heeee;
    LUT4 i30793_3_lut (.A(\mem[27] [9]), .B(\mem[26] [9]), .C(inst_reg[0]), 
         .Z(n35965)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30793_3_lut.init = 16'hcaca;
    LUT4 i30791_3_lut (.A(\mem[25] [10]), .B(\mem[24] [10]), .C(inst_reg[0]), 
         .Z(n35963)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30791_3_lut.init = 16'hcaca;
    LUT4 i30790_3_lut (.A(\mem[27] [10]), .B(\mem[26] [10]), .C(inst_reg[0]), 
         .Z(n35962)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30790_3_lut.init = 16'hcaca;
    PFUMX i30849 (.BLUT(n36019), .ALUT(n36020), .C0(inst_reg[1]), .Z(n36021));
    LUT4 i30788_3_lut (.A(\mem[25] [11]), .B(\mem[24] [11]), .C(inst_reg[0]), 
         .Z(n35960)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30788_3_lut.init = 16'hcaca;
    LUT4 i30787_3_lut (.A(\mem[27] [11]), .B(\mem[26] [11]), .C(inst_reg[0]), 
         .Z(n35959)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30787_3_lut.init = 16'hcaca;
    PFUMX i30852 (.BLUT(n36022), .ALUT(n36023), .C0(inst_reg[1]), .Z(n36024));
    LUT4 i30994_3_lut (.A(\from_fpgacfg.GPIO [0]), .B(\mem[22] [0]), .C(inst_reg[0]), 
         .Z(n36166)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30994_3_lut.init = 16'hcaca;
    LUT4 i30992_3_lut (.A(\from_fpgacfg.txant_post [0]), .B(\from_fpgacfg.txant_pre [0]), 
         .C(inst_reg[0]), .Z(n36164)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30992_3_lut.init = 16'hcaca;
    LUT4 i32301_4_lut_3_lut (.A(inst_reg[0]), .B(inst_reg[1]), .C(hw_ver_int[2]), 
         .Z(n37473)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(253[20:62])
    defparam i32301_4_lut_3_lut.init = 16'hc4c4;
    LUT4 i30991_3_lut (.A(\mem[19] [0]), .B(\mem[18] [0]), .C(inst_reg[0]), 
         .Z(n36163)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30991_3_lut.init = 16'hcaca;
    LUT4 i32297_3_lut (.A(\mem[1] [5]), .B(\mem[0] [5]), .C(inst_reg[0]), 
         .Z(n37469)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32297_3_lut.init = 16'hcaca;
    PFUMX i30861 (.BLUT(n36031), .ALUT(n36032), .C0(inst_reg[1]), .Z(n36033));
    LUT4 i32296_3_lut (.A(\mem[3] [5]), .B(\mem[2] [5]), .C(inst_reg[0]), 
         .Z(n37468)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32296_3_lut.init = 16'hcaca;
    PFUMX i30864 (.BLUT(n36034), .ALUT(n36035), .C0(inst_reg[1]), .Z(n36036));
    PFUMX i30867 (.BLUT(n36037), .ALUT(n36038), .C0(inst_reg[1]), .Z(n36039));
    LUT4 i32295_3_lut (.A(\from_fpgacfg.drct_clk_en [5]), .B(\from_fpgacfg.phase_reg_sel [5]), 
         .C(inst_reg[0]), .Z(n37467)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32295_3_lut.init = 16'hcaca;
    PFUMX i30870 (.BLUT(n36040), .ALUT(n36041), .C0(inst_reg[1]), .Z(n36042));
    PFUMX i30873 (.BLUT(n36043), .ALUT(n36044), .C0(inst_reg[1]), .Z(n36045));
    LUT4 i32294_3_lut (.A(\from_fpgacfg.ch_en [5]), .B(\from_fpgacfg.cnt_ind [0]), 
         .C(inst_reg[0]), .Z(n37466)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32294_3_lut.init = 16'hcaca;
    LUT4 i30989_3_lut (.A(\inst2_from_fpgacfg.wfm_smpl_width[0] ), .B(\from_fpgacfg.wfm_ch_en [0]), 
         .C(inst_reg[0]), .Z(n36161)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30989_3_lut.init = 16'hcaca;
    LUT4 i30988_3_lut (.A(\from_fpgacfg.sync_size [0]), .B(\mem[14] [0]), 
         .C(inst_reg[0]), .Z(n36160)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30988_3_lut.init = 16'hcaca;
    FD1P3DX din_reg__i3 (.D(din_reg[1]), .SP(REF_CLK_c_enable_1621), .CK(REF_CLK_c), 
            .CD(n41434), .Q(din_reg[2])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(133[7] 142[14])
    defparam din_reg__i3.GSR = "ENABLED";
    FD1P3DX din_reg__i4 (.D(din_reg[2]), .SP(REF_CLK_c_enable_1621), .CK(REF_CLK_c), 
            .CD(n41434), .Q(din_reg[3])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(133[7] 142[14])
    defparam din_reg__i4.GSR = "ENABLED";
    FD1P3DX din_reg__i5 (.D(din_reg[3]), .SP(REF_CLK_c_enable_1621), .CK(REF_CLK_c), 
            .CD(n41434), .Q(din_reg[4])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(133[7] 142[14])
    defparam din_reg__i5.GSR = "ENABLED";
    FD1P3DX din_reg__i6 (.D(din_reg[4]), .SP(REF_CLK_c_enable_1621), .CK(REF_CLK_c), 
            .CD(n41434), .Q(din_reg[5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(133[7] 142[14])
    defparam din_reg__i6.GSR = "ENABLED";
    FD1P3DX din_reg__i7 (.D(din_reg[5]), .SP(REF_CLK_c_enable_1621), .CK(REF_CLK_c), 
            .CD(n41434), .Q(din_reg[6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(133[7] 142[14])
    defparam din_reg__i7.GSR = "ENABLED";
    FD1P3DX din_reg__i8 (.D(din_reg[6]), .SP(REF_CLK_c_enable_1621), .CK(REF_CLK_c), 
            .CD(n41434), .Q(din_reg[7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(133[7] 142[14])
    defparam din_reg__i8.GSR = "ENABLED";
    FD1P3DX din_reg__i9 (.D(din_reg[7]), .SP(REF_CLK_c_enable_1621), .CK(REF_CLK_c), 
            .CD(n41434), .Q(din_reg[8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(133[7] 142[14])
    defparam din_reg__i9.GSR = "ENABLED";
    FD1P3DX din_reg__i10 (.D(din_reg[8]), .SP(REF_CLK_c_enable_1621), .CK(REF_CLK_c), 
            .CD(n41434), .Q(din_reg[9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(133[7] 142[14])
    defparam din_reg__i10.GSR = "ENABLED";
    FD1P3DX din_reg__i11 (.D(din_reg[9]), .SP(REF_CLK_c_enable_1621), .CK(REF_CLK_c), 
            .CD(n41434), .Q(din_reg[10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(133[7] 142[14])
    defparam din_reg__i11.GSR = "ENABLED";
    FD1P3DX din_reg__i12 (.D(din_reg[10]), .SP(REF_CLK_c_enable_1621), .CK(REF_CLK_c), 
            .CD(n41434), .Q(din_reg[11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(133[7] 142[14])
    defparam din_reg__i12.GSR = "ENABLED";
    FD1P3DX din_reg__i13 (.D(din_reg[11]), .SP(REF_CLK_c_enable_1621), .CK(REF_CLK_c), 
            .CD(n41434), .Q(din_reg[12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(133[7] 142[14])
    defparam din_reg__i13.GSR = "ENABLED";
    FD1P3DX din_reg__i14 (.D(din_reg[12]), .SP(REF_CLK_c_enable_1621), .CK(REF_CLK_c), 
            .CD(n41434), .Q(din_reg[13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(133[7] 142[14])
    defparam din_reg__i14.GSR = "ENABLED";
    FD1P3DX din_reg__i15 (.D(din_reg[13]), .SP(REF_CLK_c_enable_1621), .CK(REF_CLK_c), 
            .CD(n41434), .Q(din_reg[14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(133[7] 142[14])
    defparam din_reg__i15.GSR = "ENABLED";
    LUT4 i30986_3_lut (.A(\inst2_from_fpgacfg.smpl_nr_clr ), .B(\from_fpgacfg.smpl_width [0]), 
         .C(inst_reg[0]), .Z(n36158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30986_3_lut.init = 16'hcaca;
    LUT4 i30985_3_lut (.A(\mem[11] [0]), .B(\inst2_from_fpgacfg.rx_en ), 
         .C(inst_reg[0]), .Z(n36157)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30985_3_lut.init = 16'hcaca;
    LUT4 i30983_3_lut (.A(\from_fpgacfg.drct_clk_en [0]), .B(\from_fpgacfg.phase_reg_sel [0]), 
         .C(inst_reg[0]), .Z(n36155)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30983_3_lut.init = 16'hcaca;
    LUT4 i30982_3_lut (.A(\from_fpgacfg.ch_en [0]), .B(\from_fpgacfg.clk_ind [0]), 
         .C(inst_reg[0]), .Z(n36154)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30982_3_lut.init = 16'hcaca;
    LUT4 i30980_3_lut (.A(\mem[1] [0]), .B(\mem[0] [0]), .C(inst_reg[0]), 
         .Z(n36152)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30980_3_lut.init = 16'hcaca;
    PFUMX i30876 (.BLUT(n36046), .ALUT(n36047), .C0(inst_reg[1]), .Z(n36048));
    LUT4 i30979_3_lut (.A(\mem[3] [0]), .B(\mem[2] [0]), .C(inst_reg[0]), 
         .Z(n36151)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30979_3_lut.init = 16'hcaca;
    LUT4 mem_18__15__I_0_207_i16_2_lut (.A(\mem[18] [15]), .B(IO_0_c_0), 
         .Z(\from_fpgacfg.SPI_SS [15])) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(301[35:58])
    defparam mem_18__15__I_0_207_i16_2_lut.init = 16'hbbbb;
    LUT4 i32290_3_lut (.A(\mem[9] [5]), .B(\inst2_from_fpgacfg.mode ), .C(inst_reg[0]), 
         .Z(n37462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32290_3_lut.init = 16'hcaca;
    PFUMX i31122 (.BLUT(n36292), .ALUT(n36293), .C0(inst_reg[1]), .Z(n36294));
    PFUMX i31134 (.BLUT(n36304), .ALUT(n36305), .C0(inst_reg[1]), .Z(n36306));
    LUT4 i32289_3_lut (.A(\mem[11] [5]), .B(\mem[10] [5]), .C(inst_reg[0]), 
         .Z(n37461)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32289_3_lut.init = 16'hcaca;
    PFUMX i31137 (.BLUT(n36307), .ALUT(n36308), .C0(inst_reg[1]), .Z(n36309));
    LUT4 mem_18__15__I_0_207_i15_2_lut (.A(\mem[18] [14]), .B(IO_0_c_0), 
         .Z(\from_fpgacfg.SPI_SS [14])) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(301[35:58])
    defparam mem_18__15__I_0_207_i15_2_lut.init = 16'hbbbb;
    LUT4 i32288_3_lut (.A(\mem[13] [5]), .B(\from_fpgacfg.wfm_ch_en [5]), 
         .C(inst_reg[0]), .Z(n37460)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32288_3_lut.init = 16'hcaca;
    PFUMX i31143 (.BLUT(n36313), .ALUT(n36314), .C0(inst_reg[1]), .Z(n36315));
    LUT4 i32287_3_lut (.A(\from_fpgacfg.sync_size [5]), .B(\mem[14] [5]), 
         .C(inst_reg[0]), .Z(n37459)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32287_3_lut.init = 16'hcaca;
    LUT4 mem_18__15__I_0_207_i14_2_lut (.A(\mem[18] [13]), .B(IO_0_c_0), 
         .Z(\from_fpgacfg.SPI_SS [13])) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(301[35:58])
    defparam mem_18__15__I_0_207_i14_2_lut.init = 16'hbbbb;
    LUT4 i32283_3_lut (.A(\from_fpgacfg.txant_post [5]), .B(\from_fpgacfg.txant_pre [5]), 
         .C(inst_reg[0]), .Z(n37455)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32283_3_lut.init = 16'hcaca;
    LUT4 i32282_3_lut (.A(\inst2_from_fpgacfg.LMS1_TXEN ), .B(\mem[18] [5]), 
         .C(inst_reg[0]), .Z(n37454)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32282_3_lut.init = 16'hcaca;
    LUT4 mem_18__15__I_0_207_i13_2_lut (.A(\mem[18] [12]), .B(IO_0_c_0), 
         .Z(\from_fpgacfg.SPI_SS [12])) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(301[35:58])
    defparam mem_18__15__I_0_207_i13_2_lut.init = 16'hbbbb;
    LUT4 i32281_3_lut (.A(\mem[21] [5]), .B(\mem[20] [5]), .C(inst_reg[0]), 
         .Z(n37453)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32281_3_lut.init = 16'hcaca;
    LUT4 i32280_3_lut (.A(\from_fpgacfg.GPIO [5]), .B(\mem[22] [5]), .C(inst_reg[0]), 
         .Z(n37452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32280_3_lut.init = 16'hcaca;
    PFUMX i32074 (.BLUT(n37242), .ALUT(n37243), .C0(inst_reg[1]), .Z(n37246));
    PFUMX i32075 (.BLUT(n37244), .ALUT(n37245), .C0(inst_reg[1]), .Z(n37247));
    LUT4 mem_18__15__I_0_207_i12_2_lut (.A(\mem[18] [11]), .B(IO_0_c_0), 
         .Z(\from_fpgacfg.SPI_SS [11])) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(301[35:58])
    defparam mem_18__15__I_0_207_i12_2_lut.init = 16'hbbbb;
    PFUMX i32081 (.BLUT(n37249), .ALUT(n37250), .C0(inst_reg[1]), .Z(n37253));
    PFUMX i32082 (.BLUT(n37251), .ALUT(n37252), .C0(inst_reg[1]), .Z(n37254));
    LUT4 i32276_3_lut (.A(\mem[1] [6]), .B(\mem[0] [6]), .C(inst_reg[0]), 
         .Z(n37448)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32276_3_lut.init = 16'hcaca;
    PFUMX i32088 (.BLUT(n37256), .ALUT(n37257), .C0(inst_reg[1]), .Z(n37260));
    LUT4 i32275_3_lut (.A(\mem[3] [6]), .B(\mem[2] [6]), .C(inst_reg[0]), 
         .Z(n37447)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32275_3_lut.init = 16'hcaca;
    LUT4 i32274_3_lut (.A(\from_fpgacfg.drct_clk_en [6]), .B(\from_fpgacfg.phase_reg_sel [6]), 
         .C(inst_reg[0]), .Z(n37446)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32274_3_lut.init = 16'hcaca;
    LUT4 i32273_3_lut (.A(\from_fpgacfg.ch_en [6]), .B(\from_fpgacfg.cnt_ind [1]), 
         .C(inst_reg[0]), .Z(n37445)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32273_3_lut.init = 16'hcaca;
    LUT4 i32269_3_lut (.A(\mem[9] [6]), .B(\inst2_from_fpgacfg.ddr_en ), 
         .C(inst_reg[0]), .Z(n37441)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32269_3_lut.init = 16'hcaca;
    LUT4 i32268_3_lut (.A(\mem[11] [6]), .B(\mem[10] [6]), .C(inst_reg[0]), 
         .Z(n37440)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32268_3_lut.init = 16'hcaca;
    LUT4 i32267_3_lut (.A(\mem[13] [6]), .B(\from_fpgacfg.wfm_ch_en [6]), 
         .C(inst_reg[0]), .Z(n37439)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32267_3_lut.init = 16'hcaca;
    PFUMX i32089 (.BLUT(n37258), .ALUT(n37259), .C0(inst_reg[1]), .Z(n37261));
    LUT4 i32266_3_lut (.A(\from_fpgacfg.sync_size [6]), .B(\mem[14] [6]), 
         .C(inst_reg[0]), .Z(n37438)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32266_3_lut.init = 16'hcaca;
    PFUMX i32095 (.BLUT(n37263), .ALUT(n37264), .C0(inst_reg[1]), .Z(n37267));
    LUT4 i32262_3_lut (.A(\from_fpgacfg.txant_post [6]), .B(\from_fpgacfg.txant_pre [6]), 
         .C(inst_reg[0]), .Z(n37434)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32262_3_lut.init = 16'hcaca;
    LUT4 i32261_3_lut (.A(\inst2_from_fpgacfg.LMS1_RXEN ), .B(\mem[18] [6]), 
         .C(inst_reg[0]), .Z(n37433)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32261_3_lut.init = 16'hcaca;
    LUT4 i32260_3_lut (.A(\mem[21] [6]), .B(\mem[20] [6]), .C(inst_reg[0]), 
         .Z(n37432)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32260_3_lut.init = 16'hcaca;
    PFUMX i32096 (.BLUT(n37265), .ALUT(n37266), .C0(inst_reg[1]), .Z(n37268));
    LUT4 i32259_3_lut (.A(\from_fpgacfg.GPIO [6]), .B(\mem[22] [6]), .C(inst_reg[0]), 
         .Z(n37431)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32259_3_lut.init = 16'hcaca;
    LUT4 i32255_3_lut (.A(\mem[1] [7]), .B(\mem[0] [7]), .C(inst_reg[0]), 
         .Z(n37427)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32255_3_lut.init = 16'hcaca;
    LUT4 i32254_3_lut (.A(\mem[3] [7]), .B(\mem[2] [7]), .C(inst_reg[0]), 
         .Z(n37426)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32254_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1033 (.A(n41182), .B(inst_reg[4]), .C(n41431), 
         .D(n41443), .Z(REF_CLK_c_enable_631)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1033.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1034 (.A(n41182), .B(inst_reg[4]), .C(n41446), 
         .D(n41443), .Z(REF_CLK_c_enable_646)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1034.init = 16'h0002;
    LUT4 i1_2_lut_3_lut_4_lut_adj_1035 (.A(n41182), .B(inst_reg[4]), .C(n41447), 
         .D(n41443), .Z(REF_CLK_c_enable_661)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1035.init = 16'h0002;
    PFUMX i32102 (.BLUT(n37270), .ALUT(n37271), .C0(inst_reg[1]), .Z(n37274));
    LUT4 i1_2_lut_3_lut_4_lut_adj_1036 (.A(n41182), .B(inst_reg[4]), .C(n41384), 
         .D(n41443), .Z(REF_CLK_c_enable_676)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_1036.init = 16'h0002;
    PFUMX i32103 (.BLUT(n37272), .ALUT(n37273), .C0(inst_reg[1]), .Z(n37275));
    LUT4 i32253_3_lut (.A(\from_fpgacfg.drct_clk_en [7]), .B(\from_fpgacfg.phase_reg_sel [7]), 
         .C(inst_reg[0]), .Z(n37425)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32253_3_lut.init = 16'hcaca;
    LUT4 i32252_3_lut (.A(\from_fpgacfg.ch_en [7]), .B(\from_fpgacfg.cnt_ind [2]), 
         .C(inst_reg[0]), .Z(n37424)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32252_3_lut.init = 16'hcaca;
    PFUMX i32109 (.BLUT(n37277), .ALUT(n37278), .C0(inst_reg[1]), .Z(n37281));
    LUT4 i32248_3_lut (.A(\mem[9] [7]), .B(\inst2_from_fpgacfg.trxiq_pulse ), 
         .C(inst_reg[0]), .Z(n37420)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32248_3_lut.init = 16'hcaca;
    LUT4 i32247_3_lut (.A(\mem[11] [7]), .B(\mem[10] [7]), .C(inst_reg[0]), 
         .Z(n37419)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32247_3_lut.init = 16'hcaca;
    PFUMX i32110 (.BLUT(n37279), .ALUT(n37280), .C0(inst_reg[1]), .Z(n37282));
    PFUMX i32116 (.BLUT(n37284), .ALUT(n37285), .C0(inst_reg[1]), .Z(n37288));
    PFUMX i32117 (.BLUT(n37286), .ALUT(n37287), .C0(inst_reg[1]), .Z(n37289));
    PFUMX i32123 (.BLUT(n37291), .ALUT(n37292), .C0(inst_reg[1]), .Z(n37295));
    LUT4 i32246_3_lut (.A(\mem[13] [7]), .B(\from_fpgacfg.wfm_ch_en [7]), 
         .C(inst_reg[0]), .Z(n37418)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32246_3_lut.init = 16'hcaca;
    LUT4 i32245_3_lut (.A(\from_fpgacfg.sync_size [7]), .B(\mem[14] [7]), 
         .C(inst_reg[0]), .Z(n37417)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32245_3_lut.init = 16'hcaca;
    LUT4 i32241_3_lut (.A(\from_fpgacfg.txant_post [7]), .B(\from_fpgacfg.txant_pre [7]), 
         .C(inst_reg[0]), .Z(n37413)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32241_3_lut.init = 16'hcaca;
    LUT4 i32240_3_lut (.A(\mem[19] [7]), .B(\mem[18] [7]), .C(inst_reg[0]), 
         .Z(n37412)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32240_3_lut.init = 16'hcaca;
    PFUMX i32124 (.BLUT(n37293), .ALUT(n37294), .C0(inst_reg[1]), .Z(n37296));
    PFUMX i32130 (.BLUT(n37298), .ALUT(n37299), .C0(inst_reg[1]), .Z(n37302));
    PFUMX i32131 (.BLUT(n37300), .ALUT(n37301), .C0(inst_reg[1]), .Z(n37303));
    LUT4 i32239_3_lut (.A(\mem[21] [7]), .B(\mem[20] [7]), .C(inst_reg[0]), 
         .Z(n37411)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32239_3_lut.init = 16'hcaca;
    PFUMX i32137 (.BLUT(n37305), .ALUT(n37306), .C0(inst_reg[1]), .Z(n37309));
    LUT4 i32238_3_lut (.A(\from_fpgacfg.GPIO [7]), .B(\mem[22] [7]), .C(inst_reg[0]), 
         .Z(n37410)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32238_3_lut.init = 16'hcaca;
    LUT4 i32234_3_lut (.A(\mem[1] [8]), .B(\mem[0] [8]), .C(inst_reg[0]), 
         .Z(n37406)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32234_3_lut.init = 16'hcaca;
    LUT4 i32233_3_lut (.A(\mem[3] [8]), .B(\mem[2] [8]), .C(inst_reg[0]), 
         .Z(n37405)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32233_3_lut.init = 16'hcaca;
    LUT4 i32232_3_lut (.A(\from_fpgacfg.drct_clk_en [8]), .B(\from_fpgacfg.phase_reg_sel [8]), 
         .C(inst_reg[0]), .Z(n37404)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32232_3_lut.init = 16'hcaca;
    PFUMX i32138 (.BLUT(n37307), .ALUT(n37308), .C0(inst_reg[1]), .Z(n37310));
    LUT4 i32231_3_lut (.A(\from_fpgacfg.ch_en [8]), .B(\from_fpgacfg.cnt_ind [3]), 
         .C(inst_reg[0]), .Z(n37403)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32231_3_lut.init = 16'hcaca;
    PFUMX i32144 (.BLUT(n37312), .ALUT(n37313), .C0(inst_reg[1]), .Z(n37316));
    LUT4 i32227_3_lut (.A(\mem[9] [8]), .B(\inst2_from_fpgacfg.mimo_int_en ), 
         .C(inst_reg[0]), .Z(n37399)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32227_3_lut.init = 16'hcaca;
    LUT4 i32226_3_lut (.A(\mem[11] [8]), .B(\inst2_from_fpgacfg.rx_ptrn_en ), 
         .C(inst_reg[0]), .Z(n37398)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32226_3_lut.init = 16'hcaca;
    PFUMX i32145 (.BLUT(n37314), .ALUT(n37315), .C0(inst_reg[1]), .Z(n37317));
    LUT4 i32225_3_lut (.A(\mem[13] [8]), .B(\from_fpgacfg.wfm_ch_en [8]), 
         .C(inst_reg[0]), .Z(n37397)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32225_3_lut.init = 16'hcaca;
    PFUMX i32151 (.BLUT(n37319), .ALUT(n37320), .C0(inst_reg[1]), .Z(n37323));
    LUT4 i32224_3_lut (.A(\from_fpgacfg.sync_size [8]), .B(\mem[14] [8]), 
         .C(inst_reg[0]), .Z(n37396)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32224_3_lut.init = 16'hcaca;
    PFUMX i32152 (.BLUT(n37321), .ALUT(n37322), .C0(inst_reg[1]), .Z(n37324));
    LUT4 mem_18__15__I_0_207_i11_2_lut (.A(\mem[18] [10]), .B(IO_0_c_0), 
         .Z(\from_fpgacfg.SPI_SS [10])) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(301[35:58])
    defparam mem_18__15__I_0_207_i11_2_lut.init = 16'hbbbb;
    PFUMX i32158 (.BLUT(n37326), .ALUT(n37327), .C0(inst_reg[1]), .Z(n37330));
    LUT4 i32220_3_lut (.A(\from_fpgacfg.txant_post [8]), .B(\from_fpgacfg.txant_pre [8]), 
         .C(inst_reg[0]), .Z(n37392)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32220_3_lut.init = 16'hcaca;
    LUT4 i32219_3_lut (.A(\mem[19] [8]), .B(\mem[18] [8]), .C(inst_reg[0]), 
         .Z(n37391)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32219_3_lut.init = 16'hcaca;
    LUT4 i32218_3_lut (.A(\mem[21] [8]), .B(\mem[20] [8]), .C(inst_reg[0]), 
         .Z(n37390)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32218_3_lut.init = 16'hcaca;
    PFUMX i32159 (.BLUT(n37328), .ALUT(n37329), .C0(inst_reg[1]), .Z(n37331));
    LUT4 i32217_3_lut (.A(\from_fpgacfg.GPIO [8]), .B(\mem[22] [8]), .C(inst_reg[0]), 
         .Z(n37389)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32217_3_lut.init = 16'hcaca;
    PFUMX i32165 (.BLUT(n37333), .ALUT(n37334), .C0(inst_reg[1]), .Z(n37337));
    PFUMX i32166 (.BLUT(n37335), .ALUT(n37336), .C0(inst_reg[1]), .Z(n37338));
    PFUMX i32172 (.BLUT(n37340), .ALUT(n37341), .C0(inst_reg[1]), .Z(n37344));
    PFUMX i32173 (.BLUT(n37342), .ALUT(n37343), .C0(inst_reg[1]), .Z(n37345));
    PFUMX i32179 (.BLUT(n37347), .ALUT(n37348), .C0(inst_reg[1]), .Z(n37351));
    PFUMX i32180 (.BLUT(n37349), .ALUT(n37350), .C0(inst_reg[1]), .Z(n37352));
    PFUMX i32186 (.BLUT(n37354), .ALUT(n37355), .C0(inst_reg[1]), .Z(n37358));
    PFUMX i32187 (.BLUT(n37356), .ALUT(n37357), .C0(inst_reg[1]), .Z(n37359));
    PFUMX i32193 (.BLUT(n37361), .ALUT(n37362), .C0(inst_reg[1]), .Z(n37365));
    PFUMX i32194 (.BLUT(n37363), .ALUT(n37364), .C0(inst_reg[1]), .Z(n37366));
    PFUMX i32200 (.BLUT(n37368), .ALUT(n37369), .C0(inst_reg[1]), .Z(n37372));
    LUT4 i32026_3_lut_4_lut_else_4_lut (.A(inst_reg[1]), .B(inst_reg[2]), 
         .C(\mem[25] [3]), .D(\mem[27] [3]), .Z(n41453)) /* synthesis lut_function=(A ((C)+!B)+!A (B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam i32026_3_lut_4_lut_else_4_lut.init = 16'he6a2;
    PFUMX i32201 (.BLUT(n37370), .ALUT(n37371), .C0(inst_reg[1]), .Z(n37373));
    PFUMX i32207 (.BLUT(n37375), .ALUT(n37376), .C0(inst_reg[1]), .Z(n37379));
    PFUMX i32208 (.BLUT(n37377), .ALUT(n37378), .C0(inst_reg[1]), .Z(n37380));
    PFUMX i32214 (.BLUT(n37382), .ALUT(n37383), .C0(inst_reg[1]), .Z(n37386));
    LUT4 i14743_2_lut_rep_1026 (.A(inst_reg[0]), .B(inst_reg[1]), .Z(n41431)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14743_2_lut_rep_1026.init = 16'h8888;
    PFUMX i32215 (.BLUT(n37384), .ALUT(n37385), .C0(inst_reg[1]), .Z(n37387));
    PFUMX i32221 (.BLUT(n37389), .ALUT(n37390), .C0(inst_reg[1]), .Z(n37393));
    PFUMX i32222 (.BLUT(n37391), .ALUT(n37392), .C0(inst_reg[1]), .Z(n37394));
    PFUMX i32228 (.BLUT(n37396), .ALUT(n37397), .C0(inst_reg[1]), .Z(n37400));
    LUT4 i32033_3_lut_4_lut_then_4_lut (.A(inst_reg[1]), .B(inst_reg[2]), 
         .C(\mem[24] [1]), .D(\from_fpgacfg.FPGA_LED1_CTRL [1]), .Z(n41457)) /* synthesis lut_function=(A (B (C))+!A (B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam i32033_3_lut_4_lut_then_4_lut.init = 16'hc480;
    LUT4 i32033_3_lut_4_lut_else_4_lut (.A(inst_reg[1]), .B(inst_reg[2]), 
         .C(\mem[25] [1]), .D(\mem[27] [1]), .Z(n41456)) /* synthesis lut_function=(A ((C)+!B)+!A (B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam i32033_3_lut_4_lut_else_4_lut.init = 16'he6a2;
    PFUMX i32229 (.BLUT(n37398), .ALUT(n37399), .C0(inst_reg[1]), .Z(n37401));
    PFUMX i32235 (.BLUT(n37403), .ALUT(n37404), .C0(inst_reg[1]), .Z(n37407));
    PFUMX i32236 (.BLUT(n37405), .ALUT(n37406), .C0(inst_reg[1]), .Z(n37408));
    PFUMX i32242 (.BLUT(n37410), .ALUT(n37411), .C0(inst_reg[1]), .Z(n37414));
    LUT4 i1_2_lut_rep_1038 (.A(inst_reg[2]), .B(inst_reg[3]), .Z(n41443)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(253[20:62])
    defparam i1_2_lut_rep_1038.init = 16'heeee;
    LUT4 i1_2_lut_3_lut (.A(inst_reg[2]), .B(inst_reg[3]), .C(inst_reg[4]), 
         .Z(n31780)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(253[20:62])
    defparam i1_2_lut_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_3_lut_adj_1037 (.A(inst_reg[3]), .B(inst_reg[2]), .C(inst_reg[4]), 
         .Z(n30140)) /* synthesis lut_function=(A+!(B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(253[20:62])
    defparam i1_2_lut_3_lut_adj_1037.init = 16'hbfbf;
    LUT4 i1_2_lut_3_lut_adj_1038 (.A(inst_reg[3]), .B(inst_reg[2]), .C(inst_reg[4]), 
         .Z(n30139)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(253[20:62])
    defparam i1_2_lut_3_lut_adj_1038.init = 16'hfbfb;
    PFUMX i32243 (.BLUT(n37412), .ALUT(n37413), .C0(inst_reg[1]), .Z(n37415));
    PFUMX i32249 (.BLUT(n37417), .ALUT(n37418), .C0(inst_reg[1]), .Z(n37421));
    PFUMX i32250 (.BLUT(n37419), .ALUT(n37420), .C0(inst_reg[1]), .Z(n37422));
    PFUMX i32256 (.BLUT(n37424), .ALUT(n37425), .C0(inst_reg[1]), .Z(n37428));
    PFUMX i32257 (.BLUT(n37426), .ALUT(n37427), .C0(inst_reg[1]), .Z(n37429));
    PFUMX i32263 (.BLUT(n37431), .ALUT(n37432), .C0(inst_reg[1]), .Z(n37435));
    PFUMX i32264 (.BLUT(n37433), .ALUT(n37434), .C0(inst_reg[1]), .Z(n37436));
    PFUMX i32270 (.BLUT(n37438), .ALUT(n37439), .C0(inst_reg[1]), .Z(n37442));
    PFUMX i32271 (.BLUT(n37440), .ALUT(n37441), .C0(inst_reg[1]), .Z(n37443));
    LUT4 equal_238_i6_2_lut_rep_1041 (.A(inst_reg[0]), .B(inst_reg[1]), 
         .Z(n41446)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(253[20:62])
    defparam equal_238_i6_2_lut_rep_1041.init = 16'hbbbb;
    LUT4 i15518_2_lut_3_lut (.A(inst_reg[3]), .B(inst_reg[4]), .C(inst_reg[2]), 
         .Z(n11264)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15518_2_lut_3_lut.init = 16'h8080;
    PFUMX i32277 (.BLUT(n37445), .ALUT(n37446), .C0(inst_reg[1]), .Z(n37449));
    PFUMX i32278 (.BLUT(n37447), .ALUT(n37448), .C0(inst_reg[1]), .Z(n37450));
    LUT4 i1_2_lut_3_lut_adj_1039 (.A(inst_reg[3]), .B(inst_reg[4]), .C(inst_reg[2]), 
         .Z(n11789)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_adj_1039.init = 16'hf7f7;
    LUT4 equal_239_i6_2_lut_rep_1042 (.A(inst_reg[0]), .B(inst_reg[1]), 
         .Z(n41447)) /* synthesis lut_function=((B)+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(253[20:62])
    defparam equal_239_i6_2_lut_rep_1042.init = 16'hdddd;
    PFUMX i32284 (.BLUT(n37452), .ALUT(n37453), .C0(inst_reg[1]), .Z(n37456));
    PFUMX i32285 (.BLUT(n37454), .ALUT(n37455), .C0(inst_reg[1]), .Z(n37457));
    PFUMX i32291 (.BLUT(n37459), .ALUT(n37460), .C0(inst_reg[1]), .Z(n37463));
    PFUMX i32292 (.BLUT(n37461), .ALUT(n37462), .C0(inst_reg[1]), .Z(n37464));
    PFUMX i30981 (.BLUT(n36151), .ALUT(n36152), .C0(inst_reg[1]), .Z(n36153));
    PFUMX i30984 (.BLUT(n36154), .ALUT(n36155), .C0(inst_reg[1]), .Z(n36156));
    PFUMX i30987 (.BLUT(n36157), .ALUT(n36158), .C0(inst_reg[1]), .Z(n36159));
    LUT4 i1_2_lut_4_lut (.A(inst_reg[2]), .B(n41174), .C(inst_reg[3]), 
         .D(n41384), .Z(REF_CLK_c_enable_205)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0080;
    PFUMX i30990 (.BLUT(n36160), .ALUT(n36161), .C0(inst_reg[1]), .Z(n36162));
    LUT4 i1_2_lut_4_lut_adj_1040 (.A(inst_reg[2]), .B(n41174), .C(inst_reg[3]), 
         .D(n41431), .Z(REF_CLK_c_enable_174)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_1040.init = 16'h8000;
    LUT4 i1_2_lut_4_lut_adj_1041 (.A(inst_reg[2]), .B(n41174), .C(inst_reg[3]), 
         .D(n41446), .Z(REF_CLK_c_enable_119)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_1041.init = 16'h0080;
    LUT4 i1_2_lut_4_lut_adj_1042 (.A(inst_reg[2]), .B(n41174), .C(inst_reg[3]), 
         .D(n41447), .Z(REF_CLK_c_enable_101)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_1042.init = 16'h0080;
    PFUMX i32298 (.BLUT(n37466), .ALUT(n37467), .C0(inst_reg[1]), .Z(n37470));
    PFUMX i32299 (.BLUT(n37468), .ALUT(n37469), .C0(inst_reg[1]), .Z(n37471));
    LUT4 i32213_3_lut (.A(\mem[1] [9]), .B(\mem[0] [9]), .C(inst_reg[0]), 
         .Z(n37385)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32213_3_lut.init = 16'hcaca;
    LUT4 i32212_3_lut (.A(\mem[3] [9]), .B(\mem[2] [9]), .C(inst_reg[0]), 
         .Z(n37384)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32212_3_lut.init = 16'hcaca;
    PFUMX i30993 (.BLUT(n36163), .ALUT(n36164), .C0(inst_reg[1]), .Z(n36165));
    PFUMX i30996 (.BLUT(n36166), .ALUT(n36167), .C0(inst_reg[1]), .Z(n36168));
    LUT4 i32211_3_lut (.A(\from_fpgacfg.drct_clk_en [9]), .B(\from_fpgacfg.phase_reg_sel [9]), 
         .C(inst_reg[0]), .Z(n37383)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32211_3_lut.init = 16'hcaca;
    PFUMX i31002 (.BLUT(n36172), .ALUT(n36173), .C0(inst_reg[1]), .Z(n36174));
    LUT4 i32210_3_lut (.A(\from_fpgacfg.ch_en [9]), .B(\from_fpgacfg.cnt_ind [4]), 
         .C(inst_reg[0]), .Z(n37382)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32210_3_lut.init = 16'hcaca;
    PFUMX i32303 (.BLUT(n8), .ALUT(n9), .C0(inst_reg[1]), .Z(n37475));
    PFUMX i32304 (.BLUT(n11), .ALUT(n12), .C0(inst_reg[1]), .Z(n37476));
    LUT4 mux_16_Mux_2_i26_3_lut (.A(\mem[3] [2]), .B(\mem[2] [2]), .C(inst_reg[0]), 
         .Z(n26)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(162[13] 168[22])
    defparam mux_16_Mux_2_i26_3_lut.init = 16'hcaca;
    PFUMX i32305 (.BLUT(n16), .ALUT(n17), .C0(inst_reg[1]), .Z(n37477));
    PFUMX i32306 (.BLUT(n19), .ALUT(n20), .C0(inst_reg[1]), .Z(n37478));
    PFUMX dout_reg_15__I_0_208_i6 (.BLUT(n36049), .ALUT(dout_reg_15__N_5274[5]), 
          .C0(n37957), .Z(dout_reg_15__N_4993[5])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;
    PFUMX dout_reg_15__I_0_208_i7 (.BLUT(n36298), .ALUT(dout_reg_15__N_5274[6]), 
          .C0(n37958), .Z(dout_reg_15__N_4993[6])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;
    PFUMX dout_reg_15__I_0_208_i8 (.BLUT(n36295), .ALUT(dout_reg_15__N_5274[7]), 
          .C0(n36453), .Z(dout_reg_15__N_4993[7])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;
    PFUMX dout_reg_15__I_0_208_i9 (.BLUT(n36289), .ALUT(dout_reg_15__N_5274[8]), 
          .C0(n37958), .Z(dout_reg_15__N_4993[8])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;
    PFUMX dout_reg_15__I_0_208_i10 (.BLUT(n36286), .ALUT(dout_reg_15__N_5274[9]), 
          .C0(n37957), .Z(dout_reg_15__N_4993[9])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;
    PFUMX dout_reg_15__I_0_208_i11 (.BLUT(n36025), .ALUT(dout_reg_15__N_5274[10]), 
          .C0(n37957), .Z(dout_reg_15__N_4993[10])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;
    PFUMX dout_reg_15__I_0_208_i12 (.BLUT(n36010), .ALUT(dout_reg_15__N_5274[11]), 
          .C0(n37958), .Z(dout_reg_15__N_4993[11])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;
    PFUMX dout_reg_15__I_0_208_i13 (.BLUT(n35956), .ALUT(dout_reg_15__N_5274[12]), 
          .C0(n36453), .Z(dout_reg_15__N_4993[12])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;
    PFUMX dout_reg_15__I_0_208_i14 (.BLUT(n36310), .ALUT(dout_reg_15__N_5274[13]), 
          .C0(n36453), .Z(dout_reg_15__N_4993[13])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;
    LUT4 i32206_3_lut (.A(\mem[9] [9]), .B(\inst2_from_fpgacfg.synch_dis ), 
         .C(inst_reg[0]), .Z(n37378)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32206_3_lut.init = 16'hcaca;
    PFUMX dout_reg_15__I_0_208_i15 (.BLUT(n36301), .ALUT(dout_reg_15__N_5274[14]), 
          .C0(n37958), .Z(dout_reg_15__N_4993[14])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;
    LUT4 i32205_3_lut (.A(\mem[11] [9]), .B(\inst2_from_fpgacfg.tx_ptrn_en ), 
         .C(inst_reg[0]), .Z(n37377)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32205_3_lut.init = 16'hcaca;
    PFUMX dout_reg_15__I_0_208_i16 (.BLUT(n36274), .ALUT(dout_reg_15__N_5274[15]), 
          .C0(n37957), .Z(dout_reg_15__N_4993[15])) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=28, LSE_LLINE=110, LSE_RLINE=110 */ ;
    LUT4 i32204_3_lut (.A(\mem[13] [9]), .B(\from_fpgacfg.wfm_ch_en [9]), 
         .C(inst_reg[0]), .Z(n37376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32204_3_lut.init = 16'hcaca;
    PFUMX i32307 (.BLUT(n23), .ALUT(n24), .C0(inst_reg[1]), .Z(n37479));
    LUT4 i32203_3_lut (.A(\from_fpgacfg.sync_size [9]), .B(\mem[14] [9]), 
         .C(inst_reg[0]), .Z(n37375)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32203_3_lut.init = 16'hcaca;
    LUT4 i32199_3_lut (.A(\from_fpgacfg.txant_post [9]), .B(\from_fpgacfg.txant_pre [9]), 
         .C(inst_reg[0]), .Z(n37371)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32199_3_lut.init = 16'hcaca;
    LUT4 i32198_3_lut (.A(\mem[19] [9]), .B(\mem[18] [9]), .C(inst_reg[0]), 
         .Z(n37370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32198_3_lut.init = 16'hcaca;
    LUT4 i32197_3_lut (.A(\mem[21] [9]), .B(\mem[20] [9]), .C(inst_reg[0]), 
         .Z(n37369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32197_3_lut.init = 16'hcaca;
    LUT4 i32196_3_lut (.A(\from_fpgacfg.GPIO [9]), .B(\mem[22] [9]), .C(inst_reg[0]), 
         .Z(n37368)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32196_3_lut.init = 16'hcaca;
    LUT4 i32192_3_lut (.A(\mem[1] [10]), .B(\mem[0] [10]), .C(inst_reg[0]), 
         .Z(n37364)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i32192_3_lut.init = 16'hcaca;
    mcfg32wm_fsm fsm (.n11745(n11745), .dout_reg({dout_reg}), .dout_reg_15__N_5274({dout_reg_15__N_5274}), 
            .\dout_reg_15__N_4993[1] (dout_reg_15__N_4993[1]), .\dout_reg_15__N_4993[2] (dout_reg_15__N_4993[2]), 
            .\dout_reg_15__N_4993[3] (dout_reg_15__N_4993[3]), .\dout_reg_15__N_4993[0] (dout_reg_15__N_4993[0]), 
            .\dout_reg_15__N_4993[4] (dout_reg_15__N_4993[4]), .n36302(n36302), 
            .n36311(n36311), .REF_CLK_c(REF_CLK_c), .REF_CLK_c_enable_1453(REF_CLK_c_enable_1453), 
            .n45086(n45086), .n35957(n35957), .n36011(n36011), .n36287(n36287), 
            .n36290(n36290), .n36296(n36296), .n36299(n36299), .n36050(n36050), 
            .n36275(n36275), .n36026(n36026), .n1833(n1800[31]), .n10865(n10865), 
            .\inst_reg[11] (inst_reg[11]), .\inst_reg[13] (inst_reg[13]), 
            .\inst_reg[12] (inst_reg[12]), .\inst_reg[10] (inst_reg[10]), 
            .\inst_reg[9] (inst_reg[9]), .\inst_reg[14] (inst_reg[14]), 
            .\inst_reg[6] (inst_reg[6]), .\inst_reg[8] (inst_reg[8]), .n2023(n2023), 
            .n1848(n1800[16]), .rx_shift_data_31__N_4339(rx_shift_data_31__N_4339), 
            .\inst_reg[7] (inst_reg[7]), .\inst_reg[5] (inst_reg[5]), .n41219(n41219), 
            .IO_MISO_c(IO_MISO_c), .n45179(n45179), .\inst_reg[15] (\inst_reg[15] ), 
            .n41182(n41182), .n35448(n35448), .REF_CLK_c_enable_1621(REF_CLK_c_enable_1621), 
            .sclk_N_5010_enable_16(sclk_N_5010_enable_16), .\inst_reg[4] (inst_reg[4]), 
            .n37958(n37958), .n37957(n37957), .n36453(n36453), .USER_BUTTON_c(USER_BUTTON_c), 
            .n41434(n41434), .IO_0_c_0(IO_0_c_0));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(104[9:21])
    
endmodule
//
// Verilog Description of module mcfg32wm_fsm
//

module mcfg32wm_fsm (n11745, dout_reg, dout_reg_15__N_5274, \dout_reg_15__N_4993[1] , 
            \dout_reg_15__N_4993[2] , \dout_reg_15__N_4993[3] , \dout_reg_15__N_4993[0] , 
            \dout_reg_15__N_4993[4] , n36302, n36311, REF_CLK_c, REF_CLK_c_enable_1453, 
            n45086, n35957, n36011, n36287, n36290, n36296, n36299, 
            n36050, n36275, n36026, n1833, n10865, \inst_reg[11] , 
            \inst_reg[13] , \inst_reg[12] , \inst_reg[10] , \inst_reg[9] , 
            \inst_reg[14] , \inst_reg[6] , \inst_reg[8] , n2023, n1848, 
            rx_shift_data_31__N_4339, \inst_reg[7] , \inst_reg[5] , n41219, 
            IO_MISO_c, n45179, \inst_reg[15] , n41182, n35448, REF_CLK_c_enable_1621, 
            sclk_N_5010_enable_16, \inst_reg[4] , n37958, n37957, n36453, 
            USER_BUTTON_c, n41434, IO_0_c_0);
    output n11745;
    input [15:0]dout_reg;
    output [15:0]dout_reg_15__N_5274;
    output \dout_reg_15__N_4993[1] ;
    output \dout_reg_15__N_4993[2] ;
    output \dout_reg_15__N_4993[3] ;
    output \dout_reg_15__N_4993[0] ;
    output \dout_reg_15__N_4993[4] ;
    input n36302;
    input n36311;
    input REF_CLK_c;
    input REF_CLK_c_enable_1453;
    input n45086;
    input n35957;
    input n36011;
    input n36287;
    input n36290;
    input n36296;
    input n36299;
    input n36050;
    input n36275;
    input n36026;
    output n1833;
    output n10865;
    input \inst_reg[11] ;
    input \inst_reg[13] ;
    input \inst_reg[12] ;
    input \inst_reg[10] ;
    input \inst_reg[9] ;
    input \inst_reg[14] ;
    input \inst_reg[6] ;
    input \inst_reg[8] ;
    output n2023;
    output n1848;
    input rx_shift_data_31__N_4339;
    input \inst_reg[7] ;
    input \inst_reg[5] ;
    input n41219;
    output IO_MISO_c;
    input n45179;
    input \inst_reg[15] ;
    output n41182;
    output n35448;
    output REF_CLK_c_enable_1621;
    output sclk_N_5010_enable_16;
    input \inst_reg[4] ;
    output n37958;
    output n37957;
    output n36453;
    input USER_BUTTON_c;
    output n41434;
    input IO_0_c_0;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    
    wire n41257;
    wire [63:0]n1800;
    
    wire stateo_5__N_5806, n35392, n35406, n31594, n35390, n35402, 
        n35400, n35338, n35344, n35334, n35340, n35434, n35444, 
        n35440, n35422, n35442;
    
    LUT4 dout_reg_15__I_0_208_i2_3_lut_4_lut (.A(n11745), .B(n41257), .C(dout_reg[0]), 
         .D(dout_reg_15__N_5274[1]), .Z(\dout_reg_15__N_4993[1] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam dout_reg_15__I_0_208_i2_3_lut_4_lut.init = 16'hfd20;
    LUT4 dout_reg_15__I_0_208_i3_3_lut_4_lut (.A(n11745), .B(n41257), .C(dout_reg[1]), 
         .D(dout_reg_15__N_5274[2]), .Z(\dout_reg_15__N_4993[2] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam dout_reg_15__I_0_208_i3_3_lut_4_lut.init = 16'hfd20;
    LUT4 dout_reg_15__I_0_208_i4_3_lut_4_lut (.A(n11745), .B(n41257), .C(dout_reg[2]), 
         .D(dout_reg_15__N_5274[3]), .Z(\dout_reg_15__N_4993[3] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam dout_reg_15__I_0_208_i4_3_lut_4_lut.init = 16'hfd20;
    LUT4 dout_reg_15__I_0_208_i1_3_lut_4_lut (.A(n11745), .B(n41257), .C(dout_reg[15]), 
         .D(dout_reg_15__N_5274[0]), .Z(\dout_reg_15__N_4993[0] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam dout_reg_15__I_0_208_i1_3_lut_4_lut.init = 16'hfd20;
    LUT4 dout_reg_15__I_0_208_i5_3_lut_4_lut (.A(n11745), .B(n41257), .C(dout_reg[3]), 
         .D(dout_reg_15__N_5274[4]), .Z(\dout_reg_15__N_4993[4] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam dout_reg_15__I_0_208_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 i31131_3_lut_4_lut (.A(n11745), .B(n41257), .C(dout_reg[13]), 
         .D(n36302), .Z(dout_reg_15__N_5274[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i31131_3_lut_4_lut.init = 16'hfd20;
    LUT4 i31140_3_lut_4_lut (.A(n11745), .B(n41257), .C(dout_reg[12]), 
         .D(n36311), .Z(dout_reg_15__N_5274[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i31140_3_lut_4_lut.init = 16'hfd20;
    FD1P3BX state_FSM__i1 (.D(n45086), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .PD(stateo_5__N_5806), .Q(n1800[0]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i1.GSR = "ENABLED";
    LUT4 i30786_3_lut_4_lut (.A(n11745), .B(n41257), .C(dout_reg[11]), 
         .D(n35957), .Z(dout_reg_15__N_5274[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i30786_3_lut_4_lut.init = 16'hfd20;
    LUT4 i30840_3_lut_4_lut (.A(n11745), .B(n41257), .C(dout_reg[10]), 
         .D(n36011), .Z(dout_reg_15__N_5274[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i30840_3_lut_4_lut.init = 16'hfd20;
    LUT4 i31116_3_lut_4_lut (.A(n11745), .B(n41257), .C(dout_reg[8]), 
         .D(n36287), .Z(dout_reg_15__N_5274[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i31116_3_lut_4_lut.init = 16'hfd20;
    LUT4 i31119_3_lut_4_lut (.A(n11745), .B(n41257), .C(dout_reg[7]), 
         .D(n36290), .Z(dout_reg_15__N_5274[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i31119_3_lut_4_lut.init = 16'hfd20;
    LUT4 i31125_3_lut_4_lut (.A(n11745), .B(n41257), .C(dout_reg[6]), 
         .D(n36296), .Z(dout_reg_15__N_5274[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i31125_3_lut_4_lut.init = 16'hfd20;
    LUT4 i31128_3_lut_4_lut (.A(n11745), .B(n41257), .C(dout_reg[5]), 
         .D(n36299), .Z(dout_reg_15__N_5274[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i31128_3_lut_4_lut.init = 16'hfd20;
    LUT4 i30879_3_lut_4_lut (.A(n11745), .B(n41257), .C(dout_reg[4]), 
         .D(n36050), .Z(dout_reg_15__N_5274[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i30879_3_lut_4_lut.init = 16'hfd20;
    LUT4 i31104_3_lut_4_lut (.A(n11745), .B(n41257), .C(dout_reg[14]), 
         .D(n36275), .Z(dout_reg_15__N_5274[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i31104_3_lut_4_lut.init = 16'hfd20;
    LUT4 i30855_3_lut_4_lut (.A(n11745), .B(n41257), .C(dout_reg[9]), 
         .D(n36026), .Z(dout_reg_15__N_5274[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam i30855_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_4_lut (.A(n35392), .B(n35406), .C(n31594), .D(n35390), .Z(n11745)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(n1833), .B(n1800[26]), .Z(n35392)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_993 (.A(n1800[22]), .B(n35402), .C(n35400), .D(n1800[25]), 
         .Z(n35406)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_993.init = 16'hfffe;
    LUT4 i1_3_lut (.A(n1800[23]), .B(n1800[28]), .C(n1800[19]), .Z(n31594)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_adj_994 (.A(n1800[29]), .B(n1800[21]), .Z(n35390)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_994.init = 16'heeee;
    LUT4 i1_4_lut_adj_995 (.A(n1800[18]), .B(n1800[27]), .C(n1800[30]), 
         .D(n1800[20]), .Z(n35402)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_995.init = 16'hfffe;
    LUT4 i1_2_lut_adj_996 (.A(n1800[17]), .B(n1800[24]), .Z(n35400)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_996.init = 16'heeee;
    LUT4 i1_4_lut_adj_997 (.A(n35338), .B(n35344), .C(n35334), .D(n35340), 
         .Z(n10865)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(584[11:42])
    defparam i1_4_lut_adj_997.init = 16'hfffe;
    LUT4 i1_2_lut_adj_998 (.A(\inst_reg[11] ), .B(\inst_reg[13] ), .Z(n35338)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(584[11:42])
    defparam i1_2_lut_adj_998.init = 16'heeee;
    LUT4 i1_4_lut_adj_999 (.A(\inst_reg[12] ), .B(\inst_reg[10] ), .C(\inst_reg[9] ), 
         .D(\inst_reg[14] ), .Z(n35344)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(584[11:42])
    defparam i1_4_lut_adj_999.init = 16'hfffe;
    LUT4 i1_2_lut_adj_1000 (.A(\inst_reg[6] ), .B(\inst_reg[8] ), .Z(n35334)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(584[11:42])
    defparam i1_2_lut_adj_1000.init = 16'heeee;
    FD1P3DX state_FSM__i2 (.D(n2023), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[1]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i2.GSR = "ENABLED";
    FD1P3DX state_FSM__i3 (.D(n1800[1]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[2]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i3.GSR = "ENABLED";
    FD1P3DX state_FSM__i4 (.D(n1800[2]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[3]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i4.GSR = "ENABLED";
    FD1P3DX state_FSM__i5 (.D(n1800[3]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[4]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i5.GSR = "ENABLED";
    FD1P3DX state_FSM__i6 (.D(n1800[4]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[5]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i6.GSR = "ENABLED";
    FD1P3DX state_FSM__i7 (.D(n1800[5]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[6]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i7.GSR = "ENABLED";
    FD1P3DX state_FSM__i8 (.D(n1800[6]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[7]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i8.GSR = "ENABLED";
    FD1P3DX state_FSM__i9 (.D(n1800[7]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[8]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i9.GSR = "ENABLED";
    FD1P3DX state_FSM__i10 (.D(n1800[8]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[9]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i10.GSR = "ENABLED";
    FD1P3DX state_FSM__i11 (.D(n1800[9]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[10]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i11.GSR = "ENABLED";
    FD1P3DX state_FSM__i12 (.D(n1800[10]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[11]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i12.GSR = "ENABLED";
    FD1P3DX state_FSM__i13 (.D(n1800[11]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[12]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i13.GSR = "ENABLED";
    FD1P3DX state_FSM__i14 (.D(n1800[12]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[13]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i14.GSR = "ENABLED";
    FD1P3DX state_FSM__i15 (.D(n1800[13]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[14]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i15.GSR = "ENABLED";
    FD1P3DX state_FSM__i16 (.D(n1800[14]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[15]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i16.GSR = "ENABLED";
    FD1P3DX state_FSM__i17 (.D(n1800[15]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1848));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i17.GSR = "ENABLED";
    FD1P3DX state_FSM__i18 (.D(n1848), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[17]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i18.GSR = "ENABLED";
    FD1P3DX state_FSM__i19 (.D(n1800[17]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[18]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i19.GSR = "ENABLED";
    FD1P3DX state_FSM__i20 (.D(n1800[18]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[19]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i20.GSR = "ENABLED";
    FD1P3DX state_FSM__i21 (.D(n1800[19]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[20]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i21.GSR = "ENABLED";
    FD1P3DX state_FSM__i22 (.D(n1800[20]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[21]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i22.GSR = "ENABLED";
    FD1P3DX state_FSM__i23 (.D(n1800[21]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[22]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i23.GSR = "ENABLED";
    FD1P3DX state_FSM__i24 (.D(n1800[22]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[23]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i24.GSR = "ENABLED";
    FD1P3DX state_FSM__i25 (.D(n1800[23]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[24]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i25.GSR = "ENABLED";
    FD1P3DX state_FSM__i26 (.D(n1800[24]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[25]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i26.GSR = "ENABLED";
    FD1P3DX state_FSM__i27 (.D(n1800[25]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[26]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i27.GSR = "ENABLED";
    FD1P3DX state_FSM__i28 (.D(n1800[26]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[27]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i28.GSR = "ENABLED";
    FD1P3DX state_FSM__i29 (.D(n1800[27]), .SP(REF_CLK_c_enable_1453), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[28]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i29.GSR = "ENABLED";
    FD1P3DX state_FSM__i30 (.D(n1800[28]), .SP(rx_shift_data_31__N_4339), 
            .CK(REF_CLK_c), .CD(stateo_5__N_5806), .Q(n1800[29]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i30.GSR = "ENABLED";
    FD1P3DX state_FSM__i31 (.D(n1800[29]), .SP(rx_shift_data_31__N_4339), 
            .CK(REF_CLK_c), .CD(stateo_5__N_5806), .Q(n1800[30]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i31.GSR = "ENABLED";
    FD1P3DX state_FSM__i32 (.D(n1800[30]), .SP(rx_shift_data_31__N_4339), 
            .CK(REF_CLK_c), .CD(stateo_5__N_5806), .Q(n1833));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i32.GSR = "ENABLED";
    FD1P3DX state_FSM__i33 (.D(n1833), .SP(rx_shift_data_31__N_4339), .CK(REF_CLK_c), 
            .CD(stateo_5__N_5806), .Q(n1800[32]));   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam state_FSM__i33.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_1001 (.A(\inst_reg[7] ), .B(\inst_reg[5] ), .Z(n35340)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(584[11:42])
    defparam i1_2_lut_adj_1001.init = 16'heeee;
    LUT4 i1_4_lut_adj_1002 (.A(n41257), .B(n1800[32]), .C(dout_reg[15]), 
         .D(n41219), .Z(IO_MISO_c)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;
    defparam i1_4_lut_adj_1002.init = 16'h5040;
    LUT4 i1_2_lut_rep_777_4_lut (.A(n10865), .B(n45179), .C(\inst_reg[15] ), 
         .D(n1833), .Z(n41182)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(584[11:83])
    defparam i1_2_lut_rep_777_4_lut.init = 16'h4000;
    LUT4 i1_4_lut_adj_1003 (.A(n35434), .B(n35444), .C(n35440), .D(n35422), 
         .Z(n35448)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam i1_4_lut_adj_1003.init = 16'hfffe;
    LUT4 i1_2_lut_adj_1004 (.A(n1800[12]), .B(n1800[6]), .Z(n35434)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam i1_2_lut_adj_1004.init = 16'heeee;
    LUT4 i1_4_lut_adj_1005 (.A(n35442), .B(n1800[4]), .C(n1800[11]), .D(n1800[10]), 
         .Z(n35444)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam i1_4_lut_adj_1005.init = 16'hfffe;
    LUT4 i1_4_lut_adj_1006 (.A(n1800[3]), .B(n1800[1]), .C(n1800[2]), 
         .D(n1800[15]), .Z(n35440)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam i1_4_lut_adj_1006.init = 16'hfffe;
    LUT4 i1_2_lut_adj_1007 (.A(n1800[14]), .B(n1800[13]), .Z(n35422)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam i1_2_lut_adj_1007.init = 16'heeee;
    LUT4 i1_4_lut_adj_1008 (.A(n1800[8]), .B(n1800[7]), .C(n1800[9]), 
         .D(n1800[5]), .Z(n35442)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(92[3] 638[12])
    defparam i1_4_lut_adj_1008.init = 16'hfffe;
    LUT4 i1_2_lut_adj_1009 (.A(n1800[0]), .B(n1800[32]), .Z(n2023)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_1009.init = 16'heeee;
    LUT4 i1_2_lut_4_lut (.A(n10865), .B(n45179), .C(\inst_reg[15] ), .D(n41219), 
         .Z(REF_CLK_c_enable_1621)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/mcfg32wm_fsm.vhd(584[11:83])
    defparam i1_2_lut_4_lut.init = 16'h4000;
    LUT4 i25172_2_lut_rep_852 (.A(n10865), .B(\inst_reg[15] ), .Z(n41257)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i25172_2_lut_rep_852.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n10865), .B(\inst_reg[15] ), .C(n11745), 
         .D(n1848), .Z(sclk_N_5010_enable_16)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1110;
    LUT4 i33220_rep_194_2_lut_3_lut_4_lut (.A(n10865), .B(\inst_reg[15] ), 
         .C(\inst_reg[4] ), .D(n11745), .Z(n37958)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i33220_rep_194_2_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i33220_rep_193_2_lut_3_lut_4_lut (.A(n10865), .B(\inst_reg[15] ), 
         .C(\inst_reg[4] ), .D(n11745), .Z(n37957)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i33220_rep_193_2_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i33220_2_lut_3_lut_4_lut (.A(n10865), .B(\inst_reg[15] ), .C(\inst_reg[4] ), 
         .D(n11745), .Z(n36453)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i33220_2_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 lreset_I_0_1_lut_rep_1029 (.A(USER_BUTTON_c), .Z(n41434)) /* synthesis lut_function=(!(A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(89[10:22])
    defparam lreset_I_0_1_lut_rep_1029.init = 16'h5555;
    LUT4 sen_I_0_175_2_lut_2_lut (.A(USER_BUTTON_c), .B(IO_0_c_0), .Z(stateo_5__N_5806)) /* synthesis lut_function=((B)+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(89[10:22])
    defparam sen_I_0_175_2_lut_2_lut.init = 16'hdddd;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module platform1_vhd
//

module platform1_vhd (\SHAREDBUS_ADR_I[7] , n3, \SHAREDBUS_ADR_I[10] , 
            n41347, n41303, REF_CLK_c, REF_CLK_c_enable_1606, n41434, 
            inst1_FIFOof_wr, n41301, n41310, inst3_Full, inst1_FIFOif_rd, 
            n35647, inst3_Empty, n41298, n41300, n29, n41263, \SHAREDBUS_ADR_I[29] , 
            \SHAREDBUS_ADR_I[23] , n45101, \counter[2] , n12428, n41346, 
            n2, \selected[0] , n32312, \SHAREDBUS_ADR_I[5] , n34966, 
            n34926, \SHAREDBUS_ADR_I[22] , n34242, n41344, n41299, 
            n30231, PIO_DATAI, sclk_N_5010, IO_SCK_c, rx_shift_data_31__N_4339, 
            n41328, REF_CLK_c_enable_1453, IO_MISO_c, IO_0_c_0, GND_net, 
            VCC_net, IO_MOSI_c, n41329, n41330, n41331, n41332, 
            n41333, n41334, n41335, \SHAREDBUS_DAT_I[8] , \SHAREDBUS_DAT_I[9] , 
            \SHAREDBUS_DAT_I[10] , \SHAREDBUS_DAT_I[11] , \SHAREDBUS_DAT_I[12] , 
            \SHAREDBUS_DAT_I[13] , \SHAREDBUS_DAT_I[14] , \SHAREDBUS_DAT_I[15] , 
            n41336, n41337, n41338, n41339, n41340, n41341, n41342, 
            n41343, \SHAREDBUS_DAT_I[24] , \SHAREDBUS_DAT_I[25] , \SHAREDBUS_DAT_I[26] , 
            \SHAREDBUS_DAT_I[27] , \SHAREDBUS_DAT_I[28] , \SHAREDBUS_DAT_I[29] , 
            \SHAREDBUS_DAT_I[30] , \SHAREDBUS_DAT_I[31] , n45179, n41380, 
            \inst_reg[15] , n10865, n41191, \genblk1.read_address[10] , 
            \genblk1.write_address[10] , n3700, n5386, n5085, n3432, 
            \genblk1.state[2] , \genblk1.pmi_address[3] , \genblk1.pmi_address[4] , 
            \genblk1.pmi_address[5] , \genblk1.pmi_address[6] , \genblk1.pmi_address[7] , 
            \genblk1.pmi_address[8] , \genblk1.pmi_address[9] , \genblk1.pmi_address[10] , 
            \genblk1.pmi_address[11] , \genblk1.pmi_address[12] , \genblk1.pmi_address[13] , 
            \genblk1.pmi_address[14] , n41321, n20000, n6038, n11843, 
            n3485, n6034, n41292, n19822, n41390, n3486, n82_adj_343, 
            n45076, n8, LM32D_CYC_O, locked_N_493, \LM32D_CTI_O[0] , 
            \LM32I_ADR_O[12] , n29830, \next_cycle_type[2] , write_idx_w, 
            n41352, n41351, w_result, n41350, dcache_refill_request, 
            \operand_1_x[1] , dc_re, n41430, n41432, REF_CLK_c_enable_176, 
            n7611, n41405, REF_CLK_c_enable_164, n41356, n41355, n41353, 
            n41358, n41359, \operand_m[10] , \operand_m[9] , \operand_m[5] , 
            dcache_select_x, n41354, bie, n31279, \adder_result_x[16] , 
            \adder_result_x[17] , \adder_result_x[18] , \adder_result_x[19] , 
            \adder_result_x[20] , \adder_result_x[21] , \adder_result_x[22] , 
            \adder_result_x[23] , \adder_result_x[24] , \adder_result_x[25] , 
            \adder_result_x[26] , \adder_result_x[27] , \adder_result_x[28] , 
            \adder_result_x[29] , \adder_result_x[30] , \adder_result_x[31] , 
            n6518, n6648, branch_target_d, direction_m, n45103, n45099, 
            n41394, n41401, bie_N_3274, pc_f, n41325, n17816, n41379, 
            \shifter_result_m[21] , n41357, \left_shift_result[21] , \left_shift_result[10] , 
            b, \p[0] , \p[1] , \p[2] , \p[3] , \p[4] , \p[5] , 
            \p[6] , \p[7] , \p[8] , \p[9] , \p[10] , \p[11] , \p[12] , 
            \p[13] , \p[14] , \p[15] , \p[16] , \p[17] , \p[18] , 
            \p[19] , \p[20] , \p[21] , \p[22] , \p[23] , \p[24] , 
            \p[25] , \p[26] , \p[27] , \p[28] , \p[29] , \p[30] , 
            \a[31] , t, n38965, \d_adr_o_31__N_2278[5] , \d_adr_o_31__N_2278[9] , 
            \d_adr_o_31__N_2278[10] , \LM32D_ADR_O[17] , \LM32D_ADR_O[19] , 
            \state[0] , \state[2] , flush_set, flush_set_8__N_2513, 
            \dcache_refill_address[5] , \dcache_refill_address[9] , \dcache_refill_address[10] , 
            \tmem_write_address[1] , \tmem_write_address[5] , \tmem_write_address[6] , 
            \dmem_write_address[3] , \dmem_write_address[7] , \dmem_write_address[8] , 
            n36337, n6781, n6764, n6749, pc_d, n6760, n45105, 
            n6589, n6584, n37179, n6439, n6434, n37177, n6599, 
            n6594, n37180, n6629, n6624, n37183, n6579, n6574, 
            n37178, n6429, n6424, n37176, n6609, n6604, n37181, 
            n6619, n6614, n37182, n37185, n37184, n37188, n37187, 
            n37186, n37189, n7603, n7571, n7607, n7575, n7606, 
            n7574, n7604, n7572, n7605, n7573, n7608, n7576, n7602, 
            n7570, n7601, n7569, n7600, n7568, n7599, n7567, n7598, 
            n7566, n7597, n7565, n7596, n7564, n7595, n7563, n7594, 
            n7562, n7593, n7561, n7592, n7560, n7584, n7552, n7583, 
            n7551, n7582, n7550, n7581, n7549, n7580, n7548, n7579, 
            n7547, n7578, n7546, n7577, n7545, n6750, n7591, n7559, 
            n7590, n7558, n7589, n7557, n7588, n7556, n7587, n7555, 
            n7586, n7554, n7585, n7553, n37501, n37500, n37502, 
            n37499, n37498, n37497, n37496, n6751, n6752, n6753, 
            n6754, n6755, n6756, n6757, n6758, n6759, n6761, n6762, 
            n6763, n37495, n7672, n7640, n7673, n7641, n34_adj_327, 
            n7674, n7642, n7675, n7643, n7676, n7644, n7671, n7639, 
            n7670, n7638, n7669, n7637, n7668, n7636, n7667, n7635, 
            n7666, n7634, n7665, n7633, n7664, n7632, n7663, n7631, 
            n7662, n7630, n7661, n7629, n7660, n7628, n36, n7652, 
            n7620, n7651, n7619, n7650, n7618, n7649, n7617, n37_adj_328, 
            n7648, n7616, n7647, n7615, n7646, n7614, n7645, n7613, 
            n7659, n7627, n7658, n7626, n7657, n7625, n7656, n7624, 
            n7655, n7623, n7654, n7622, n7653, n7621, n37504, 
            n37503, n37507, n37506, n37505, n37508, n45106, \LM32I_ADR_O[17] , 
            \LM32I_ADR_O[19] , flush_set_adj_344, flush_set_8__N_1953, 
            n157, n36336, n10589, n10585, n10591, n10593, n10587, 
            n10595, n10452, LED_R_c_0, n36338, LED_G_c_0, LED_B_c_0, 
            n36339, n36340, n35006, inst1_FIFOfifo_rst, inst3_Q);
    output \SHAREDBUS_ADR_I[7] ;
    output n3;
    output \SHAREDBUS_ADR_I[10] ;
    output n41347;
    output n41303;
    input REF_CLK_c;
    output REF_CLK_c_enable_1606;
    input n41434;
    output inst1_FIFOof_wr;
    output n41301;
    output n41310;
    input inst3_Full;
    output inst1_FIFOif_rd;
    input n35647;
    input inst3_Empty;
    output n41298;
    output n41300;
    input n29;
    input n41263;
    output \SHAREDBUS_ADR_I[29] ;
    output \SHAREDBUS_ADR_I[23] ;
    output n45101;
    output \counter[2] ;
    input n12428;
    output n41346;
    output n2;
    output \selected[0] ;
    input n32312;
    output \SHAREDBUS_ADR_I[5] ;
    output n34966;
    output n34926;
    output \SHAREDBUS_ADR_I[22] ;
    input n34242;
    output n41344;
    output n41299;
    output n30231;
    output [0:0]PIO_DATAI;
    output sclk_N_5010;
    output IO_SCK_c;
    output rx_shift_data_31__N_4339;
    output n41328;
    output REF_CLK_c_enable_1453;
    input IO_MISO_c;
    output IO_0_c_0;
    input GND_net;
    input VCC_net;
    output IO_MOSI_c;
    output n41329;
    output n41330;
    output n41331;
    output n41332;
    output n41333;
    output n41334;
    output n41335;
    output \SHAREDBUS_DAT_I[8] ;
    output \SHAREDBUS_DAT_I[9] ;
    output \SHAREDBUS_DAT_I[10] ;
    output \SHAREDBUS_DAT_I[11] ;
    output \SHAREDBUS_DAT_I[12] ;
    output \SHAREDBUS_DAT_I[13] ;
    output \SHAREDBUS_DAT_I[14] ;
    output \SHAREDBUS_DAT_I[15] ;
    output n41336;
    output n41337;
    output n41338;
    output n41339;
    output n41340;
    output n41341;
    output n41342;
    output n41343;
    output \SHAREDBUS_DAT_I[24] ;
    output \SHAREDBUS_DAT_I[25] ;
    output \SHAREDBUS_DAT_I[26] ;
    output \SHAREDBUS_DAT_I[27] ;
    output \SHAREDBUS_DAT_I[28] ;
    output \SHAREDBUS_DAT_I[29] ;
    output \SHAREDBUS_DAT_I[30] ;
    output \SHAREDBUS_DAT_I[31] ;
    output n45179;
    output n41380;
    input \inst_reg[15] ;
    input n10865;
    output n41191;
    input \genblk1.read_address[10] ;
    input \genblk1.write_address[10] ;
    output n3700;
    output n5386;
    output n5085;
    output n3432;
    output \genblk1.state[2] ;
    output \genblk1.pmi_address[3] ;
    output \genblk1.pmi_address[4] ;
    output \genblk1.pmi_address[5] ;
    output \genblk1.pmi_address[6] ;
    output \genblk1.pmi_address[7] ;
    output \genblk1.pmi_address[8] ;
    output \genblk1.pmi_address[9] ;
    output \genblk1.pmi_address[10] ;
    output \genblk1.pmi_address[11] ;
    output \genblk1.pmi_address[12] ;
    output \genblk1.pmi_address[13] ;
    output \genblk1.pmi_address[14] ;
    output n41321;
    output n20000;
    output n6038;
    output n11843;
    output n3485;
    output n6034;
    output n41292;
    output n19822;
    output n41390;
    output n3486;
    input [14:0]n82_adj_343;
    output n45076;
    output n8;
    output LM32D_CYC_O;
    output locked_N_493;
    output \LM32D_CTI_O[0] ;
    output \LM32I_ADR_O[12] ;
    output n29830;
    output \next_cycle_type[2] ;
    output [4:0]write_idx_w;
    output n41352;
    output n41351;
    output [31:0]w_result;
    output n41350;
    output dcache_refill_request;
    output \operand_1_x[1] ;
    output dc_re;
    output n41430;
    input n41432;
    output REF_CLK_c_enable_176;
    output n7611;
    input n41405;
    output REF_CLK_c_enable_164;
    output n41356;
    output n41355;
    output n41353;
    output n41358;
    output n41359;
    output \operand_m[10] ;
    output \operand_m[9] ;
    output \operand_m[5] ;
    input dcache_select_x;
    output n41354;
    output bie;
    output n31279;
    output \adder_result_x[16] ;
    output \adder_result_x[17] ;
    output \adder_result_x[18] ;
    output \adder_result_x[19] ;
    output \adder_result_x[20] ;
    output \adder_result_x[21] ;
    output \adder_result_x[22] ;
    output \adder_result_x[23] ;
    output \adder_result_x[24] ;
    output \adder_result_x[25] ;
    output \adder_result_x[26] ;
    output \adder_result_x[27] ;
    output \adder_result_x[28] ;
    output \adder_result_x[29] ;
    output \adder_result_x[30] ;
    output \adder_result_x[31] ;
    input n6518;
    input n6648;
    input [31:2]branch_target_d;
    output direction_m;
    output n45103;
    output n45099;
    output n41394;
    output n41401;
    output bie_N_3274;
    output [31:2]pc_f;
    output n41325;
    input n17816;
    output n41379;
    input \shifter_result_m[21] ;
    output n41357;
    output \left_shift_result[21] ;
    output \left_shift_result[10] ;
    output [31:0]b;
    output \p[0] ;
    output \p[1] ;
    output \p[2] ;
    output \p[3] ;
    output \p[4] ;
    output \p[5] ;
    output \p[6] ;
    output \p[7] ;
    output \p[8] ;
    output \p[9] ;
    output \p[10] ;
    output \p[11] ;
    output \p[12] ;
    output \p[13] ;
    output \p[14] ;
    output \p[15] ;
    output \p[16] ;
    output \p[17] ;
    output \p[18] ;
    output \p[19] ;
    output \p[20] ;
    output \p[21] ;
    output \p[22] ;
    output \p[23] ;
    output \p[24] ;
    output \p[25] ;
    output \p[26] ;
    output \p[27] ;
    output \p[28] ;
    output \p[29] ;
    output \p[30] ;
    output \a[31] ;
    input [32:0]t;
    input n38965;
    input \d_adr_o_31__N_2278[5] ;
    input \d_adr_o_31__N_2278[9] ;
    input \d_adr_o_31__N_2278[10] ;
    output \LM32D_ADR_O[17] ;
    output \LM32D_ADR_O[19] ;
    output \state[0] ;
    output \state[2] ;
    output [8:0]flush_set;
    input [8:0]flush_set_8__N_2513;
    output \dcache_refill_address[5] ;
    output \dcache_refill_address[9] ;
    output \dcache_refill_address[10] ;
    input \tmem_write_address[1] ;
    input \tmem_write_address[5] ;
    input \tmem_write_address[6] ;
    input \dmem_write_address[3] ;
    input \dmem_write_address[7] ;
    input \dmem_write_address[8] ;
    input n36337;
    output n6781;
    output n6764;
    output n6749;
    output [31:2]pc_d;
    output n6760;
    output n45105;
    input n6589;
    input n6584;
    output n37179;
    input n6439;
    input n6434;
    output n37177;
    input n6599;
    input n6594;
    output n37180;
    input n6629;
    input n6624;
    output n37183;
    input n6579;
    input n6574;
    output n37178;
    input n6429;
    input n6424;
    output n37176;
    input n6609;
    input n6604;
    output n37181;
    input n6619;
    input n6614;
    output n37182;
    input n37185;
    input n37184;
    output n37188;
    input n37187;
    input n37186;
    output n37189;
    input n7603;
    input n7571;
    input n7607;
    input n7575;
    input n7606;
    input n7574;
    input n7604;
    input n7572;
    input n7605;
    input n7573;
    input n7608;
    input n7576;
    input n7602;
    input n7570;
    input n7601;
    input n7569;
    input n7600;
    input n7568;
    input n7599;
    input n7567;
    input n7598;
    input n7566;
    input n7597;
    input n7565;
    input n7596;
    input n7564;
    input n7595;
    input n7563;
    input n7594;
    input n7562;
    input n7593;
    input n7561;
    input n7592;
    input n7560;
    input n7584;
    input n7552;
    input n7583;
    input n7551;
    input n7582;
    input n7550;
    input n7581;
    input n7549;
    input n7580;
    input n7548;
    input n7579;
    input n7547;
    input n7578;
    input n7546;
    input n7577;
    input n7545;
    output n6750;
    input n7591;
    input n7559;
    input n7590;
    input n7558;
    input n7589;
    input n7557;
    input n7588;
    input n7556;
    input n7587;
    input n7555;
    input n7586;
    input n7554;
    input n7585;
    input n7553;
    output n37501;
    output n37500;
    output n37502;
    output n37499;
    output n37498;
    output n37497;
    output n37496;
    output n6751;
    output n6752;
    output n6753;
    output n6754;
    output n6755;
    output n6756;
    output n6757;
    output n6758;
    output n6759;
    output n6761;
    output n6762;
    output n6763;
    output n37495;
    input n7672;
    input n7640;
    input n7673;
    input n7641;
    output n34_adj_327;
    input n7674;
    input n7642;
    input n7675;
    input n7643;
    input n7676;
    input n7644;
    input n7671;
    input n7639;
    input n7670;
    input n7638;
    input n7669;
    input n7637;
    input n7668;
    input n7636;
    input n7667;
    input n7635;
    input n7666;
    input n7634;
    input n7665;
    input n7633;
    input n7664;
    input n7632;
    input n7663;
    input n7631;
    input n7662;
    input n7630;
    input n7661;
    input n7629;
    input n7660;
    input n7628;
    output n36;
    input n7652;
    input n7620;
    input n7651;
    input n7619;
    input n7650;
    input n7618;
    input n7649;
    input n7617;
    output n37_adj_328;
    input n7648;
    input n7616;
    input n7647;
    input n7615;
    input n7646;
    input n7614;
    input n7645;
    input n7613;
    input n7659;
    input n7627;
    input n7658;
    input n7626;
    input n7657;
    input n7625;
    input n7656;
    input n7624;
    input n7655;
    input n7623;
    input n7654;
    input n7622;
    input n7653;
    input n7621;
    input n37504;
    input n37503;
    output n37507;
    input n37506;
    input n37505;
    output n37508;
    output n45106;
    output \LM32I_ADR_O[17] ;
    output \LM32I_ADR_O[19] ;
    output [8:0]flush_set_adj_344;
    input [8:0]flush_set_8__N_1953;
    input [29:0]n157;
    input n36336;
    output n10589;
    output n10585;
    output n10591;
    output n10593;
    output n10587;
    output n10595;
    output n10452;
    output LED_R_c_0;
    input n36338;
    output LED_G_c_0;
    output LED_B_c_0;
    input n36339;
    input n36340;
    output n35006;
    output inst1_FIFOfifo_rst;
    input [31:0]inst3_Q;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire sclk_N_5010 /* synthesis is_inv_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(57[11:19])
    wire IO_SCK_c /* synthesis is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(28[3:9])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    
    platform1 lm32_inst (.\SHAREDBUS_ADR_I[7] (\SHAREDBUS_ADR_I[7] ), .n3(n3), 
            .\SHAREDBUS_ADR_I[10] (\SHAREDBUS_ADR_I[10] ), .n41347(n41347), 
            .n41303(n41303), .REF_CLK_c(REF_CLK_c), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .n41434(n41434), .inst1_FIFOof_wr(inst1_FIFOof_wr), .n41301(n41301), 
            .n41310(n41310), .inst3_Full(inst3_Full), .inst1_FIFOif_rd(inst1_FIFOif_rd), 
            .n35647(n35647), .inst3_Empty(inst3_Empty), .n41298(n41298), 
            .n41300(n41300), .n29(n29), .n41263(n41263), .\SHAREDBUS_ADR_I[29] (\SHAREDBUS_ADR_I[29] ), 
            .\SHAREDBUS_ADR_I[23] (\SHAREDBUS_ADR_I[23] ), .n45101(n45101), 
            .\counter[2] (\counter[2] ), .n12428(n12428), .n41346(n41346), 
            .n2(n2), .selected({Open_0, \selected[0] }), .n32312(n32312), 
            .\SHAREDBUS_ADR_I[5] (\SHAREDBUS_ADR_I[5] ), .n34966(n34966), 
            .n34926(n34926), .\SHAREDBUS_ADR_I[22] (\SHAREDBUS_ADR_I[22] ), 
            .n34242(n34242), .n41344(n41344), .n41299(n41299), .n30231(n30231), 
            .PIO_DATAI({PIO_DATAI}), .sclk_N_5010(sclk_N_5010), .IO_SCK_c(IO_SCK_c), 
            .rx_shift_data_31__N_4339(rx_shift_data_31__N_4339), .n41328(n41328), 
            .REF_CLK_c_enable_1453(REF_CLK_c_enable_1453), .IO_MISO_c(IO_MISO_c), 
            .IO_0_c_0(IO_0_c_0), .GND_net(GND_net), .VCC_net(VCC_net), 
            .IO_MOSI_c(IO_MOSI_c), .n41329(n41329), .n41330(n41330), .n41331(n41331), 
            .n41332(n41332), .n41333(n41333), .n41334(n41334), .n41335(n41335), 
            .\SHAREDBUS_DAT_I[8] (\SHAREDBUS_DAT_I[8] ), .\SHAREDBUS_DAT_I[9] (\SHAREDBUS_DAT_I[9] ), 
            .\SHAREDBUS_DAT_I[10] (\SHAREDBUS_DAT_I[10] ), .\SHAREDBUS_DAT_I[11] (\SHAREDBUS_DAT_I[11] ), 
            .\SHAREDBUS_DAT_I[12] (\SHAREDBUS_DAT_I[12] ), .\SHAREDBUS_DAT_I[13] (\SHAREDBUS_DAT_I[13] ), 
            .\SHAREDBUS_DAT_I[14] (\SHAREDBUS_DAT_I[14] ), .\SHAREDBUS_DAT_I[15] (\SHAREDBUS_DAT_I[15] ), 
            .n41336(n41336), .n41337(n41337), .n41338(n41338), .n41339(n41339), 
            .n41340(n41340), .n41341(n41341), .n41342(n41342), .n41343(n41343), 
            .\SHAREDBUS_DAT_I[24] (\SHAREDBUS_DAT_I[24] ), .\SHAREDBUS_DAT_I[25] (\SHAREDBUS_DAT_I[25] ), 
            .\SHAREDBUS_DAT_I[26] (\SHAREDBUS_DAT_I[26] ), .\SHAREDBUS_DAT_I[27] (\SHAREDBUS_DAT_I[27] ), 
            .\SHAREDBUS_DAT_I[28] (\SHAREDBUS_DAT_I[28] ), .\SHAREDBUS_DAT_I[29] (\SHAREDBUS_DAT_I[29] ), 
            .\SHAREDBUS_DAT_I[30] (\SHAREDBUS_DAT_I[30] ), .\SHAREDBUS_DAT_I[31] (\SHAREDBUS_DAT_I[31] ), 
            .n45179(n45179), .n41380(n41380), .\inst_reg[15] (\inst_reg[15] ), 
            .n10865(n10865), .n41191(n41191), .\genblk1.read_address[10] (\genblk1.read_address[10] ), 
            .\genblk1.write_address[10] (\genblk1.write_address[10] ), .n3700(n3700), 
            .n5386(n5386), .n5085(n5085), .n3432(n3432), .\genblk1.state[2] (\genblk1.state[2] ), 
            .\genblk1.pmi_address[3] (\genblk1.pmi_address[3] ), .\genblk1.pmi_address[4] (\genblk1.pmi_address[4] ), 
            .\genblk1.pmi_address[5] (\genblk1.pmi_address[5] ), .\genblk1.pmi_address[6] (\genblk1.pmi_address[6] ), 
            .\genblk1.pmi_address[7] (\genblk1.pmi_address[7] ), .\genblk1.pmi_address[8] (\genblk1.pmi_address[8] ), 
            .\genblk1.pmi_address[9] (\genblk1.pmi_address[9] ), .\genblk1.pmi_address[10] (\genblk1.pmi_address[10] ), 
            .\genblk1.pmi_address[11] (\genblk1.pmi_address[11] ), .\genblk1.pmi_address[12] (\genblk1.pmi_address[12] ), 
            .\genblk1.pmi_address[13] (\genblk1.pmi_address[13] ), .\genblk1.pmi_address[14] (\genblk1.pmi_address[14] ), 
            .n41321(n41321), .n20000(n20000), .n6038(n6038), .n11843(n11843), 
            .n3485(n3485), .n6034(n6034), .n41292(n41292), .n19822(n19822), 
            .n41390(n41390), .n3486(n3486), .n82_adj_325({n82_adj_343}), 
            .n45076(n45076), .n8(n8), .LM32D_CYC_O(LM32D_CYC_O), .locked_N_493(locked_N_493), 
            .\LM32D_CTI_O[0] (\LM32D_CTI_O[0] ), .\LM32I_ADR_O[12] (\LM32I_ADR_O[12] ), 
            .n29830(n29830), .\next_cycle_type[2] (\next_cycle_type[2] ), 
            .write_idx_w({write_idx_w}), .n41352(n41352), .n41351(n41351), 
            .w_result({w_result}), .n41350(n41350), .dcache_refill_request(dcache_refill_request), 
            .\operand_1_x[1] (\operand_1_x[1] ), .dc_re(dc_re), .n41430(n41430), 
            .n41432(n41432), .REF_CLK_c_enable_176(REF_CLK_c_enable_176), 
            .n7611(n7611), .n41405(n41405), .REF_CLK_c_enable_164(REF_CLK_c_enable_164), 
            .n41356(n41356), .n41355(n41355), .n41353(n41353), .n41358(n41358), 
            .n41359(n41359), .\operand_m[10] (\operand_m[10] ), .\operand_m[9] (\operand_m[9] ), 
            .\operand_m[5] (\operand_m[5] ), .dcache_select_x(dcache_select_x), 
            .n41354(n41354), .bie(bie), .n31279(n31279), .\adder_result_x[16] (\adder_result_x[16] ), 
            .\adder_result_x[17] (\adder_result_x[17] ), .\adder_result_x[18] (\adder_result_x[18] ), 
            .\adder_result_x[19] (\adder_result_x[19] ), .\adder_result_x[20] (\adder_result_x[20] ), 
            .\adder_result_x[21] (\adder_result_x[21] ), .\adder_result_x[22] (\adder_result_x[22] ), 
            .\adder_result_x[23] (\adder_result_x[23] ), .\adder_result_x[24] (\adder_result_x[24] ), 
            .\adder_result_x[25] (\adder_result_x[25] ), .\adder_result_x[26] (\adder_result_x[26] ), 
            .\adder_result_x[27] (\adder_result_x[27] ), .\adder_result_x[28] (\adder_result_x[28] ), 
            .\adder_result_x[29] (\adder_result_x[29] ), .\adder_result_x[30] (\adder_result_x[30] ), 
            .\adder_result_x[31] (\adder_result_x[31] ), .n6518(n6518), 
            .n6648(n6648), .branch_target_d({branch_target_d}), .direction_m(direction_m), 
            .n45103(n45103), .n45099(n45099), .n41394(n41394), .n41401(n41401), 
            .bie_N_3274(bie_N_3274), .pc_f({pc_f}), .n41325(n41325), .n17816(n17816), 
            .n41379(n41379), .\shifter_result_m[21] (\shifter_result_m[21] ), 
            .n41357(n41357), .\left_shift_result[21] (\left_shift_result[21] ), 
            .\left_shift_result[10] (\left_shift_result[10] ), .b({b}), 
            .\p[0] (\p[0] ), .\p[1] (\p[1] ), .\p[2] (\p[2] ), .\p[3] (\p[3] ), 
            .\p[4] (\p[4] ), .\p[5] (\p[5] ), .\p[6] (\p[6] ), .\p[7] (\p[7] ), 
            .\p[8] (\p[8] ), .\p[9] (\p[9] ), .\p[10] (\p[10] ), .\p[11] (\p[11] ), 
            .\p[12] (\p[12] ), .\p[13] (\p[13] ), .\p[14] (\p[14] ), .\p[15] (\p[15] ), 
            .\p[16] (\p[16] ), .\p[17] (\p[17] ), .\p[18] (\p[18] ), .\p[19] (\p[19] ), 
            .\p[20] (\p[20] ), .\p[21] (\p[21] ), .\p[22] (\p[22] ), .\p[23] (\p[23] ), 
            .\p[24] (\p[24] ), .\p[25] (\p[25] ), .\p[26] (\p[26] ), .\p[27] (\p[27] ), 
            .\p[28] (\p[28] ), .\p[29] (\p[29] ), .\p[30] (\p[30] ), .\a[31] (\a[31] ), 
            .t({t}), .n38965(n38965), .\d_adr_o_31__N_2278[5] (\d_adr_o_31__N_2278[5] ), 
            .\d_adr_o_31__N_2278[9] (\d_adr_o_31__N_2278[9] ), .\d_adr_o_31__N_2278[10] (\d_adr_o_31__N_2278[10] ), 
            .\LM32D_ADR_O[17] (\LM32D_ADR_O[17] ), .\LM32D_ADR_O[19] (\LM32D_ADR_O[19] ), 
            .\state[0] (\state[0] ), .\state[2] (\state[2] ), .flush_set({flush_set}), 
            .flush_set_8__N_2513({flush_set_8__N_2513}), .\dcache_refill_address[5] (\dcache_refill_address[5] ), 
            .\dcache_refill_address[9] (\dcache_refill_address[9] ), .\dcache_refill_address[10] (\dcache_refill_address[10] ), 
            .\tmem_write_address[1] (\tmem_write_address[1] ), .\tmem_write_address[5] (\tmem_write_address[5] ), 
            .\tmem_write_address[6] (\tmem_write_address[6] ), .\dmem_write_address[3] (\dmem_write_address[3] ), 
            .\dmem_write_address[7] (\dmem_write_address[7] ), .\dmem_write_address[8] (\dmem_write_address[8] ), 
            .n36337(n36337), .n6781(n6781), .n6764(n6764), .n6749(n6749), 
            .pc_d({pc_d}), .n6760(n6760), .n45105(n45105), .n6589(n6589), 
            .n6584(n6584), .n37179(n37179), .n6439(n6439), .n6434(n6434), 
            .n37177(n37177), .n6599(n6599), .n6594(n6594), .n37180(n37180), 
            .n6629(n6629), .n6624(n6624), .n37183(n37183), .n6579(n6579), 
            .n6574(n6574), .n37178(n37178), .n6429(n6429), .n6424(n6424), 
            .n37176(n37176), .n6609(n6609), .n6604(n6604), .n37181(n37181), 
            .n6619(n6619), .n6614(n6614), .n37182(n37182), .n37185(n37185), 
            .n37184(n37184), .n37188(n37188), .n37187(n37187), .n37186(n37186), 
            .n37189(n37189), .n7603(n7603), .n7571(n7571), .n7607(n7607), 
            .n7575(n7575), .n7606(n7606), .n7574(n7574), .n7604(n7604), 
            .n7572(n7572), .n7605(n7605), .n7573(n7573), .n7608(n7608), 
            .n7576(n7576), .n7602(n7602), .n7570(n7570), .n7601(n7601), 
            .n7569(n7569), .n7600(n7600), .n7568(n7568), .n7599(n7599), 
            .n7567(n7567), .n7598(n7598), .n7566(n7566), .n7597(n7597), 
            .n7565(n7565), .n7596(n7596), .n7564(n7564), .n7595(n7595), 
            .n7563(n7563), .n7594(n7594), .n7562(n7562), .n7593(n7593), 
            .n7561(n7561), .n7592(n7592), .n7560(n7560), .n7584(n7584), 
            .n7552(n7552), .n7583(n7583), .n7551(n7551), .n7582(n7582), 
            .n7550(n7550), .n7581(n7581), .n7549(n7549), .n7580(n7580), 
            .n7548(n7548), .n7579(n7579), .n7547(n7547), .n7578(n7578), 
            .n7546(n7546), .n7577(n7577), .n7545(n7545), .n6750(n6750), 
            .n7591(n7591), .n7559(n7559), .n7590(n7590), .n7558(n7558), 
            .n7589(n7589), .n7557(n7557), .n7588(n7588), .n7556(n7556), 
            .n7587(n7587), .n7555(n7555), .n7586(n7586), .n7554(n7554), 
            .n7585(n7585), .n7553(n7553), .n37501(n37501), .n37500(n37500), 
            .n37502(n37502), .n37499(n37499), .n37498(n37498), .n37497(n37497), 
            .n37496(n37496), .n6751(n6751), .n6752(n6752), .n6753(n6753), 
            .n6754(n6754), .n6755(n6755), .n6756(n6756), .n6757(n6757), 
            .n6758(n6758), .n6759(n6759), .n6761(n6761), .n6762(n6762), 
            .n6763(n6763), .n37495(n37495), .n7672(n7672), .n7640(n7640), 
            .n7673(n7673), .n7641(n7641), .n34_adj_309(n34_adj_327), .n7674(n7674), 
            .n7642(n7642), .n7675(n7675), .n7643(n7643), .n7676(n7676), 
            .n7644(n7644), .n7671(n7671), .n7639(n7639), .n7670(n7670), 
            .n7638(n7638), .n7669(n7669), .n7637(n7637), .n7668(n7668), 
            .n7636(n7636), .n7667(n7667), .n7635(n7635), .n7666(n7666), 
            .n7634(n7634), .n7665(n7665), .n7633(n7633), .n7664(n7664), 
            .n7632(n7632), .n7663(n7663), .n7631(n7631), .n7662(n7662), 
            .n7630(n7630), .n7661(n7661), .n7629(n7629), .n7660(n7660), 
            .n7628(n7628), .n36(n36), .n7652(n7652), .n7620(n7620), 
            .n7651(n7651), .n7619(n7619), .n7650(n7650), .n7618(n7618), 
            .n7649(n7649), .n7617(n7617), .n37_adj_310(n37_adj_328), .n7648(n7648), 
            .n7616(n7616), .n7647(n7647), .n7615(n7615), .n7646(n7646), 
            .n7614(n7614), .n7645(n7645), .n7613(n7613), .n7659(n7659), 
            .n7627(n7627), .n7658(n7658), .n7626(n7626), .n7657(n7657), 
            .n7625(n7625), .n7656(n7656), .n7624(n7624), .n7655(n7655), 
            .n7623(n7623), .n7654(n7654), .n7622(n7622), .n7653(n7653), 
            .n7621(n7621), .n37504(n37504), .n37503(n37503), .n37507(n37507), 
            .n37506(n37506), .n37505(n37505), .n37508(n37508), .n45106(n45106), 
            .\LM32I_ADR_O[17] (\LM32I_ADR_O[17] ), .\LM32I_ADR_O[19] (\LM32I_ADR_O[19] ), 
            .flush_set_adj_326({flush_set_adj_344}), .flush_set_8__N_1953({flush_set_8__N_1953}), 
            .n157({n157}), .n36336(n36336), .n10589(n10589), .n10585(n10585), 
            .n10591(n10591), .n10593(n10593), .n10587(n10587), .n10595(n10595), 
            .n10452(n10452), .LED_R_c_0(LED_R_c_0), .n36338(n36338), .LED_G_c_0(LED_G_c_0), 
            .LED_B_c_0(LED_B_c_0), .n36339(n36339), .n36340(n36340), .n35006(n35006), 
            .inst1_FIFOfifo_rst(inst1_FIFOfifo_rst), .inst3_Q({inst3_Q})) /* synthesis syn_module_defined=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1_vhd.vhd(54[13:22])
    
endmodule
//
// Verilog Description of module platform1
//

module platform1 (\SHAREDBUS_ADR_I[7] , n3, \SHAREDBUS_ADR_I[10] , n41347, 
            n41303, REF_CLK_c, REF_CLK_c_enable_1606, n41434, inst1_FIFOof_wr, 
            n41301, n41310, inst3_Full, inst1_FIFOif_rd, n35647, inst3_Empty, 
            n41298, n41300, n29, n41263, \SHAREDBUS_ADR_I[29] , \SHAREDBUS_ADR_I[23] , 
            n45101, \counter[2] , n12428, n41346, n2, selected, 
            n32312, \SHAREDBUS_ADR_I[5] , n34966, n34926, \SHAREDBUS_ADR_I[22] , 
            n34242, n41344, n41299, n30231, PIO_DATAI, sclk_N_5010, 
            IO_SCK_c, rx_shift_data_31__N_4339, n41328, REF_CLK_c_enable_1453, 
            IO_MISO_c, IO_0_c_0, GND_net, VCC_net, IO_MOSI_c, n41329, 
            n41330, n41331, n41332, n41333, n41334, n41335, \SHAREDBUS_DAT_I[8] , 
            \SHAREDBUS_DAT_I[9] , \SHAREDBUS_DAT_I[10] , \SHAREDBUS_DAT_I[11] , 
            \SHAREDBUS_DAT_I[12] , \SHAREDBUS_DAT_I[13] , \SHAREDBUS_DAT_I[14] , 
            \SHAREDBUS_DAT_I[15] , n41336, n41337, n41338, n41339, 
            n41340, n41341, n41342, n41343, \SHAREDBUS_DAT_I[24] , 
            \SHAREDBUS_DAT_I[25] , \SHAREDBUS_DAT_I[26] , \SHAREDBUS_DAT_I[27] , 
            \SHAREDBUS_DAT_I[28] , \SHAREDBUS_DAT_I[29] , \SHAREDBUS_DAT_I[30] , 
            \SHAREDBUS_DAT_I[31] , n45179, n41380, \inst_reg[15] , n10865, 
            n41191, \genblk1.read_address[10] , \genblk1.write_address[10] , 
            n3700, n5386, n5085, n3432, \genblk1.state[2] , \genblk1.pmi_address[3] , 
            \genblk1.pmi_address[4] , \genblk1.pmi_address[5] , \genblk1.pmi_address[6] , 
            \genblk1.pmi_address[7] , \genblk1.pmi_address[8] , \genblk1.pmi_address[9] , 
            \genblk1.pmi_address[10] , \genblk1.pmi_address[11] , \genblk1.pmi_address[12] , 
            \genblk1.pmi_address[13] , \genblk1.pmi_address[14] , n41321, 
            n20000, n6038, n11843, n3485, n6034, n41292, n19822, 
            n41390, n3486, n82_adj_325, n45076, n8, LM32D_CYC_O, 
            locked_N_493, \LM32D_CTI_O[0] , \LM32I_ADR_O[12] , n29830, 
            \next_cycle_type[2] , write_idx_w, n41352, n41351, w_result, 
            n41350, dcache_refill_request, \operand_1_x[1] , dc_re, 
            n41430, n41432, REF_CLK_c_enable_176, n7611, n41405, REF_CLK_c_enable_164, 
            n41356, n41355, n41353, n41358, n41359, \operand_m[10] , 
            \operand_m[9] , \operand_m[5] , dcache_select_x, n41354, 
            bie, n31279, \adder_result_x[16] , \adder_result_x[17] , 
            \adder_result_x[18] , \adder_result_x[19] , \adder_result_x[20] , 
            \adder_result_x[21] , \adder_result_x[22] , \adder_result_x[23] , 
            \adder_result_x[24] , \adder_result_x[25] , \adder_result_x[26] , 
            \adder_result_x[27] , \adder_result_x[28] , \adder_result_x[29] , 
            \adder_result_x[30] , \adder_result_x[31] , n6518, n6648, 
            branch_target_d, direction_m, n45103, n45099, n41394, 
            n41401, bie_N_3274, pc_f, n41325, n17816, n41379, \shifter_result_m[21] , 
            n41357, \left_shift_result[21] , \left_shift_result[10] , 
            b, \p[0] , \p[1] , \p[2] , \p[3] , \p[4] , \p[5] , 
            \p[6] , \p[7] , \p[8] , \p[9] , \p[10] , \p[11] , \p[12] , 
            \p[13] , \p[14] , \p[15] , \p[16] , \p[17] , \p[18] , 
            \p[19] , \p[20] , \p[21] , \p[22] , \p[23] , \p[24] , 
            \p[25] , \p[26] , \p[27] , \p[28] , \p[29] , \p[30] , 
            \a[31] , t, n38965, \d_adr_o_31__N_2278[5] , \d_adr_o_31__N_2278[9] , 
            \d_adr_o_31__N_2278[10] , \LM32D_ADR_O[17] , \LM32D_ADR_O[19] , 
            \state[0] , \state[2] , flush_set, flush_set_8__N_2513, 
            \dcache_refill_address[5] , \dcache_refill_address[9] , \dcache_refill_address[10] , 
            \tmem_write_address[1] , \tmem_write_address[5] , \tmem_write_address[6] , 
            \dmem_write_address[3] , \dmem_write_address[7] , \dmem_write_address[8] , 
            n36337, n6781, n6764, n6749, pc_d, n6760, n45105, 
            n6589, n6584, n37179, n6439, n6434, n37177, n6599, 
            n6594, n37180, n6629, n6624, n37183, n6579, n6574, 
            n37178, n6429, n6424, n37176, n6609, n6604, n37181, 
            n6619, n6614, n37182, n37185, n37184, n37188, n37187, 
            n37186, n37189, n7603, n7571, n7607, n7575, n7606, 
            n7574, n7604, n7572, n7605, n7573, n7608, n7576, n7602, 
            n7570, n7601, n7569, n7600, n7568, n7599, n7567, n7598, 
            n7566, n7597, n7565, n7596, n7564, n7595, n7563, n7594, 
            n7562, n7593, n7561, n7592, n7560, n7584, n7552, n7583, 
            n7551, n7582, n7550, n7581, n7549, n7580, n7548, n7579, 
            n7547, n7578, n7546, n7577, n7545, n6750, n7591, n7559, 
            n7590, n7558, n7589, n7557, n7588, n7556, n7587, n7555, 
            n7586, n7554, n7585, n7553, n37501, n37500, n37502, 
            n37499, n37498, n37497, n37496, n6751, n6752, n6753, 
            n6754, n6755, n6756, n6757, n6758, n6759, n6761, n6762, 
            n6763, n37495, n7672, n7640, n7673, n7641, n34_adj_309, 
            n7674, n7642, n7675, n7643, n7676, n7644, n7671, n7639, 
            n7670, n7638, n7669, n7637, n7668, n7636, n7667, n7635, 
            n7666, n7634, n7665, n7633, n7664, n7632, n7663, n7631, 
            n7662, n7630, n7661, n7629, n7660, n7628, n36, n7652, 
            n7620, n7651, n7619, n7650, n7618, n7649, n7617, n37_adj_310, 
            n7648, n7616, n7647, n7615, n7646, n7614, n7645, n7613, 
            n7659, n7627, n7658, n7626, n7657, n7625, n7656, n7624, 
            n7655, n7623, n7654, n7622, n7653, n7621, n37504, 
            n37503, n37507, n37506, n37505, n37508, n45106, \LM32I_ADR_O[17] , 
            \LM32I_ADR_O[19] , flush_set_adj_326, flush_set_8__N_1953, 
            n157, n36336, n10589, n10585, n10591, n10593, n10587, 
            n10595, n10452, LED_R_c_0, n36338, LED_G_c_0, LED_B_c_0, 
            n36339, n36340, n35006, inst1_FIFOfifo_rst, inst3_Q) /* synthesis syn_module_defined=1 */ ;
    output \SHAREDBUS_ADR_I[7] ;
    output n3;
    output \SHAREDBUS_ADR_I[10] ;
    output n41347;
    output n41303;
    input REF_CLK_c;
    output REF_CLK_c_enable_1606;
    input n41434;
    output inst1_FIFOof_wr;
    output n41301;
    output n41310;
    input inst3_Full;
    output inst1_FIFOif_rd;
    input n35647;
    input inst3_Empty;
    output n41298;
    output n41300;
    input n29;
    input n41263;
    output \SHAREDBUS_ADR_I[29] ;
    output \SHAREDBUS_ADR_I[23] ;
    output n45101;
    output \counter[2] ;
    input n12428;
    output n41346;
    output n2;
    output [1:0]selected;
    input n32312;
    output \SHAREDBUS_ADR_I[5] ;
    output n34966;
    output n34926;
    output \SHAREDBUS_ADR_I[22] ;
    input n34242;
    output n41344;
    output n41299;
    output n30231;
    output [0:0]PIO_DATAI;
    output sclk_N_5010;
    output IO_SCK_c;
    output rx_shift_data_31__N_4339;
    output n41328;
    output REF_CLK_c_enable_1453;
    input IO_MISO_c;
    output IO_0_c_0;
    input GND_net;
    input VCC_net;
    output IO_MOSI_c;
    output n41329;
    output n41330;
    output n41331;
    output n41332;
    output n41333;
    output n41334;
    output n41335;
    output \SHAREDBUS_DAT_I[8] ;
    output \SHAREDBUS_DAT_I[9] ;
    output \SHAREDBUS_DAT_I[10] ;
    output \SHAREDBUS_DAT_I[11] ;
    output \SHAREDBUS_DAT_I[12] ;
    output \SHAREDBUS_DAT_I[13] ;
    output \SHAREDBUS_DAT_I[14] ;
    output \SHAREDBUS_DAT_I[15] ;
    output n41336;
    output n41337;
    output n41338;
    output n41339;
    output n41340;
    output n41341;
    output n41342;
    output n41343;
    output \SHAREDBUS_DAT_I[24] ;
    output \SHAREDBUS_DAT_I[25] ;
    output \SHAREDBUS_DAT_I[26] ;
    output \SHAREDBUS_DAT_I[27] ;
    output \SHAREDBUS_DAT_I[28] ;
    output \SHAREDBUS_DAT_I[29] ;
    output \SHAREDBUS_DAT_I[30] ;
    output \SHAREDBUS_DAT_I[31] ;
    output n45179;
    output n41380;
    input \inst_reg[15] ;
    input n10865;
    output n41191;
    input \genblk1.read_address[10] ;
    input \genblk1.write_address[10] ;
    output n3700;
    output n5386;
    output n5085;
    output n3432;
    output \genblk1.state[2] ;
    output \genblk1.pmi_address[3] ;
    output \genblk1.pmi_address[4] ;
    output \genblk1.pmi_address[5] ;
    output \genblk1.pmi_address[6] ;
    output \genblk1.pmi_address[7] ;
    output \genblk1.pmi_address[8] ;
    output \genblk1.pmi_address[9] ;
    output \genblk1.pmi_address[10] ;
    output \genblk1.pmi_address[11] ;
    output \genblk1.pmi_address[12] ;
    output \genblk1.pmi_address[13] ;
    output \genblk1.pmi_address[14] ;
    output n41321;
    output n20000;
    output n6038;
    output n11843;
    output n3485;
    output n6034;
    output n41292;
    output n19822;
    output n41390;
    output n3486;
    input [14:0]n82_adj_325;
    output n45076;
    output n8;
    output LM32D_CYC_O;
    output locked_N_493;
    output \LM32D_CTI_O[0] ;
    output \LM32I_ADR_O[12] ;
    output n29830;
    output \next_cycle_type[2] ;
    output [4:0]write_idx_w;
    output n41352;
    output n41351;
    output [31:0]w_result;
    output n41350;
    output dcache_refill_request;
    output \operand_1_x[1] ;
    output dc_re;
    output n41430;
    input n41432;
    output REF_CLK_c_enable_176;
    output n7611;
    input n41405;
    output REF_CLK_c_enable_164;
    output n41356;
    output n41355;
    output n41353;
    output n41358;
    output n41359;
    output \operand_m[10] ;
    output \operand_m[9] ;
    output \operand_m[5] ;
    input dcache_select_x;
    output n41354;
    output bie;
    output n31279;
    output \adder_result_x[16] ;
    output \adder_result_x[17] ;
    output \adder_result_x[18] ;
    output \adder_result_x[19] ;
    output \adder_result_x[20] ;
    output \adder_result_x[21] ;
    output \adder_result_x[22] ;
    output \adder_result_x[23] ;
    output \adder_result_x[24] ;
    output \adder_result_x[25] ;
    output \adder_result_x[26] ;
    output \adder_result_x[27] ;
    output \adder_result_x[28] ;
    output \adder_result_x[29] ;
    output \adder_result_x[30] ;
    output \adder_result_x[31] ;
    input n6518;
    input n6648;
    input [31:2]branch_target_d;
    output direction_m;
    output n45103;
    output n45099;
    output n41394;
    output n41401;
    output bie_N_3274;
    output [31:2]pc_f;
    output n41325;
    input n17816;
    output n41379;
    input \shifter_result_m[21] ;
    output n41357;
    output \left_shift_result[21] ;
    output \left_shift_result[10] ;
    output [31:0]b;
    output \p[0] ;
    output \p[1] ;
    output \p[2] ;
    output \p[3] ;
    output \p[4] ;
    output \p[5] ;
    output \p[6] ;
    output \p[7] ;
    output \p[8] ;
    output \p[9] ;
    output \p[10] ;
    output \p[11] ;
    output \p[12] ;
    output \p[13] ;
    output \p[14] ;
    output \p[15] ;
    output \p[16] ;
    output \p[17] ;
    output \p[18] ;
    output \p[19] ;
    output \p[20] ;
    output \p[21] ;
    output \p[22] ;
    output \p[23] ;
    output \p[24] ;
    output \p[25] ;
    output \p[26] ;
    output \p[27] ;
    output \p[28] ;
    output \p[29] ;
    output \p[30] ;
    output \a[31] ;
    input [32:0]t;
    input n38965;
    input \d_adr_o_31__N_2278[5] ;
    input \d_adr_o_31__N_2278[9] ;
    input \d_adr_o_31__N_2278[10] ;
    output \LM32D_ADR_O[17] ;
    output \LM32D_ADR_O[19] ;
    output \state[0] ;
    output \state[2] ;
    output [8:0]flush_set;
    input [8:0]flush_set_8__N_2513;
    output \dcache_refill_address[5] ;
    output \dcache_refill_address[9] ;
    output \dcache_refill_address[10] ;
    input \tmem_write_address[1] ;
    input \tmem_write_address[5] ;
    input \tmem_write_address[6] ;
    input \dmem_write_address[3] ;
    input \dmem_write_address[7] ;
    input \dmem_write_address[8] ;
    input n36337;
    output n6781;
    output n6764;
    output n6749;
    output [31:2]pc_d;
    output n6760;
    output n45105;
    input n6589;
    input n6584;
    output n37179;
    input n6439;
    input n6434;
    output n37177;
    input n6599;
    input n6594;
    output n37180;
    input n6629;
    input n6624;
    output n37183;
    input n6579;
    input n6574;
    output n37178;
    input n6429;
    input n6424;
    output n37176;
    input n6609;
    input n6604;
    output n37181;
    input n6619;
    input n6614;
    output n37182;
    input n37185;
    input n37184;
    output n37188;
    input n37187;
    input n37186;
    output n37189;
    input n7603;
    input n7571;
    input n7607;
    input n7575;
    input n7606;
    input n7574;
    input n7604;
    input n7572;
    input n7605;
    input n7573;
    input n7608;
    input n7576;
    input n7602;
    input n7570;
    input n7601;
    input n7569;
    input n7600;
    input n7568;
    input n7599;
    input n7567;
    input n7598;
    input n7566;
    input n7597;
    input n7565;
    input n7596;
    input n7564;
    input n7595;
    input n7563;
    input n7594;
    input n7562;
    input n7593;
    input n7561;
    input n7592;
    input n7560;
    input n7584;
    input n7552;
    input n7583;
    input n7551;
    input n7582;
    input n7550;
    input n7581;
    input n7549;
    input n7580;
    input n7548;
    input n7579;
    input n7547;
    input n7578;
    input n7546;
    input n7577;
    input n7545;
    output n6750;
    input n7591;
    input n7559;
    input n7590;
    input n7558;
    input n7589;
    input n7557;
    input n7588;
    input n7556;
    input n7587;
    input n7555;
    input n7586;
    input n7554;
    input n7585;
    input n7553;
    output n37501;
    output n37500;
    output n37502;
    output n37499;
    output n37498;
    output n37497;
    output n37496;
    output n6751;
    output n6752;
    output n6753;
    output n6754;
    output n6755;
    output n6756;
    output n6757;
    output n6758;
    output n6759;
    output n6761;
    output n6762;
    output n6763;
    output n37495;
    input n7672;
    input n7640;
    input n7673;
    input n7641;
    output n34_adj_309;
    input n7674;
    input n7642;
    input n7675;
    input n7643;
    input n7676;
    input n7644;
    input n7671;
    input n7639;
    input n7670;
    input n7638;
    input n7669;
    input n7637;
    input n7668;
    input n7636;
    input n7667;
    input n7635;
    input n7666;
    input n7634;
    input n7665;
    input n7633;
    input n7664;
    input n7632;
    input n7663;
    input n7631;
    input n7662;
    input n7630;
    input n7661;
    input n7629;
    input n7660;
    input n7628;
    output n36;
    input n7652;
    input n7620;
    input n7651;
    input n7619;
    input n7650;
    input n7618;
    input n7649;
    input n7617;
    output n37_adj_310;
    input n7648;
    input n7616;
    input n7647;
    input n7615;
    input n7646;
    input n7614;
    input n7645;
    input n7613;
    input n7659;
    input n7627;
    input n7658;
    input n7626;
    input n7657;
    input n7625;
    input n7656;
    input n7624;
    input n7655;
    input n7623;
    input n7654;
    input n7622;
    input n7653;
    input n7621;
    input n37504;
    input n37503;
    output n37507;
    input n37506;
    input n37505;
    output n37508;
    output n45106;
    output \LM32I_ADR_O[17] ;
    output \LM32I_ADR_O[19] ;
    output [8:0]flush_set_adj_326;
    input [8:0]flush_set_8__N_1953;
    input [29:0]n157;
    input n36336;
    output n10589;
    output n10585;
    output n10591;
    output n10593;
    output n10587;
    output n10595;
    output n10452;
    output LED_R_c_0;
    input n36338;
    output LED_G_c_0;
    output LED_B_c_0;
    input n36339;
    input n36340;
    output n35006;
    output inst1_FIFOfifo_rst;
    input [31:0]inst3_Q;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire sclk_N_5010 /* synthesis is_inv_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(57[11:19])
    wire IO_SCK_c /* synthesis is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(28[3:9])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    wire [31:0]ebrEBR_DAT_O;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(417[13:25])
    wire [31:0]\genblk1.write_data_d ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(241[43:55])
    
    wire \genblk1.raw_hazard , n9, n11, n32332, n41210, n41186, 
        n36988;
    wire [31:0]\genblk1.read_data ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(245[31:40])
    
    wire n36343;
    wire [2:0]n1;
    
    wire n41276, n41253, n32798, n35761, n35868, n41234;
    wire [31:0]SHAREDBUS_ADR_I;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(361[13:28])
    
    wire n37927, n37931, n37930, n37929, n37928, n41189, n37926, 
        n37932, n41251, n33368, n41273, n41269, n41277, n41242, 
        n35840, n35712, n15, n35890, n41246, n41279, n34698, n9_adj_6341;
    wire [31:0]\genblk1.EBR_DAT_I_d ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(248[31:42])
    wire [3:0]\genblk1.EBR_SEL_I_d ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(249[16:27])
    wire [7:0]\genblk1.write_data_23__N_3549 ;
    
    wire n41236, n33088;
    wire [31:0]n4865;
    
    wire n32980, n32940, n33100, n33060, n32864, n33020, n11_adj_6342, 
        n9_adj_6343, n9_adj_6344, n34704, n35633, n34702, n19, n34692, 
        n41237, n41278, n34672, n31779, n34664, n35908, n34650, 
        n41225, n35796, n41272, n41274, n34632, fiford_reg, n11769, 
        n19808, n41194, n37907, n37909, n35942, n31833, n61, n31955, 
        n35844, n35888, n41259, n35886, n32728, n32900, n41262, 
        n32898, n30762, n32882, n41265, n32890, n41264, n32200, 
        n32194, REF_CLK_c_enable_424, n41268, n32192, n41267, n32174, 
        n37910, n37911, n37908, n37912, n37913, n41235, n32028, 
        n32032, n35186, n35808, n41492, n41493, n41220, n32694, 
        n32690, n35912, n32464, n41193, n41195;
    wire [31:0]n1030;
    
    wire ebrEBR_ACK_O;
    wire [31:0]n1063;
    
    wire n21, n16, n34992, PIO_DATAI_0__N_3822;
    wire [7:0]\genblk1.write_data_15__N_3565 ;
    
    wire n11_adj_6346, spiSPI_ACK_O, n32084, n47;
    wire [31:0]n997;
    wire [31:0]n1096;
    
    wire n41181;
    wire [31:0]SHAREDBUS_ACK_O_N_91;
    wire [31:0]spiSPI_DAT_O;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(440[13:25])
    
    wire FIFOwb_en;
    wire [31:0]FIFOwb_DAT_O;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(451[13:25])
    
    wire n3_adj_6347, n34304;
    wire [31:0]reg_00;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(80[15:21])
    
    wire n41185, n34226, n15_adj_6348, n3_adj_6349, n34302, n15_adj_6350, 
        n3_adj_6351, n34378, n15_adj_6352, n3_adj_6353, n34416, n15_adj_6354, 
        n9_adj_6355, n3_adj_6356, n34340, n15_adj_6357, n3_adj_6358, 
        n34264, n15_adj_6359, n33030, n17, n33366, n13, n3_adj_6360, 
        n34036, n15_adj_6361, n3_adj_6362, n34188, n15_adj_6363, n32874, 
        n23, n33070, n17_adj_6364, n33252, n13_adj_6365, n33110, 
        n17_adj_6366, n33290, n13_adj_6367, n32950, n17_adj_6368, 
        n33404, n13_adj_6369, n30944, n6;
    wire [7:0]GPOout_pins;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1_vhd.vhd(11[3:14])
    
    wire n34150, n4, n30948, n6_adj_6370, n34454, n4_adj_6371, n32990, 
        n15_adj_6372, n33328, n11_adj_6373, n30951, n6_adj_6374, n34074, 
        n4_adj_6375, n30949, n6_adj_6376, n33998, n4_adj_6377;
    wire [31:0]n295;
    
    wire n11_adj_6378, n17_adj_6379, n17_adj_6380, n17_adj_6381, n17_adj_6382, 
        n17_adj_6383, n15_adj_6384, n17_adj_6385, n17_adj_6386, n17_adj_6387, 
        n17_adj_6388, n17_adj_6389, n14, n17_adj_6390, n14_adj_6391, 
        n26, n11_adj_6392, n17_adj_6393, n14_adj_6394, n9_adj_6395, 
        n5, n11_adj_6396, n17_adj_6397, n14_adj_6398, n11_adj_6399, 
        n11_adj_6400;
    wire [7:0]\genblk1.write_data_31__N_3533 ;
    wire [0:0]n949;
    
    wire n30241, n31750, n13990;
    wire [31:0]LM32D_ADR_O;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(389[13:24])
    
    wire n5_adj_6401, n11_adj_6402, n9_adj_6403, n22, n9_adj_6404, 
        n22_adj_6405, n9_adj_6406;
    wire [31:0]LM32I_ADR_O;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(376[13:24])
    
    wire n22_adj_6407, n9_adj_6408, n2_adj_6409, n11_adj_6410, n2_adj_6411, 
        n11_adj_6412, n22_adj_6413, n9_adj_6414, n5_adj_6415, n11_adj_6416, 
        n2_adj_6417, n11_adj_6418, n26_adj_6419, n11_adj_6420, n2_adj_6421, 
        n11_adj_6422;
    wire [31:0]n361;
    
    wire n11_adj_6423, n5_adj_6424, n11_adj_6425, n11_adj_6426, n25, 
        n11_adj_6427, n5_adj_6428, n11_adj_6429, n11_adj_6430, n25_adj_6431, 
        n11_adj_6432, n25_adj_6433, n11_adj_6434, n5_adj_6435, n11_adj_6436, 
        n25_adj_6437, n11_adj_6438, n25_adj_6439, n11_adj_6440, n22_adj_6441, 
        n11_adj_6442, n32038, n32036, n30986, n25_adj_6443, n11_adj_6444, 
        n9_adj_6445, n11_adj_6446, n35200, n35892, n31476, n35184, 
        n41270, n41266, n41254, n11_adj_6447, n9_adj_6448, n9_adj_6449, 
        n7, n9_adj_6450, n11_adj_6451, n9_adj_6452, n35605, n35649, 
        n35160, write_ack_N_4649, n41260, n35136, n35236, fiford, 
        n35222, n35204;
    wire [0:0]n954;
    
    wire GPIOGPIO_ACK_O, n41252, n34960, n41275, n41239, n31, n13_adj_6453, 
        n32326, n34372, n32322, n32304, n32318, n32788, n35884, 
        n32774, n33846, n35739, read_ack, n41180, write_ack, n36351, 
        n34104, n34444, n34112, n34078, n34396, n34236;
    wire [31:0]reg_04;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(81[15:21])
    
    wire n33990, n33964, n34066, n34040, n35910, n34446, n34420, 
        n34142, n34116, n35724, n41304, n41345, n34816, n33864, 
        n35577, n35854, n33954, n31183, n33332, n33356, n32814, 
        n32828, n8_c;
    wire [31:0]SHAREDBUS_DAT_O;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(363[13:28])
    
    wire n8_adj_6454, n8_adj_6455, n8_adj_6456, n8_adj_6457, n8_adj_6458, 
        n8_adj_6459, n8_adj_6460, n8_adj_6461, n8_adj_6462, n8_adj_6463, 
        n8_adj_6464, n8_adj_6465, n8_adj_6466, n8_adj_6467, n8_adj_6468, 
        n8_adj_6469, n8_adj_6470, n3_adj_6471, n8_adj_6472, n8_adj_6473, 
        n3_adj_6474, n3_adj_6475, n3_adj_6476, n8_adj_6477, n33214, 
        n3_adj_6478, n8_adj_6479, n3_adj_6480, n8_adj_6481, n3_adj_6482, 
        n3_adj_6483, n11_adj_6484, n14_adj_6485, n13_adj_6486, n19_adj_6487, 
        n13_adj_6488, n19_adj_6489, n13_adj_6490, n19_adj_6491, n13_adj_6492, 
        n19_adj_6493, n33948, n11_adj_6494, n17_adj_6495, n13_adj_6496, 
        n19_adj_6497, n13_adj_6498, n19_adj_6499, n13_adj_6500, n19_adj_6501, 
        n13_adj_6502, n19_adj_6503, n9_adj_6504, n19_adj_6505;
    wire [31:0]GPOwb_DAT_O;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(432[13:24])
    wire [31:0]n328;
    
    wire n8_adj_6506, n8_adj_6507, n17_adj_6508, n8_adj_6509, n8_adj_6510, 
        n19_adj_6511, n19_adj_6512, n19_adj_6513, n16_adj_6514, n16_adj_6515, 
        n19_adj_6516, n16_adj_6517, n16_adj_6518, n34180, n34154, 
        n16_adj_6519, n16_adj_6520, n16_adj_6521, n16_adj_6522, n34028, 
        n34002, n34256, n34230, n34332, n34306, n34408, n34382, 
        n34370, n34344, n34294, n34268, n34218, n34192, n32074, 
        n35930, n32054, n35866, write_ack_adj_6523, read_ack_adj_6524, 
        dw10_cs_N_4471, dw00_cs_N_4467, n30156, n35042, n34742, SPI_INT_O_N_4422, 
        SPI_INT_O_N_4417, SPI_INT_O_N_4421;
    wire [0:0]n953;
    
    wire \genblk1.wait_one_tick_done ;
    wire [7:0]\genblk1.write_data_7__N_3573 ;
    
    wire n41324, n41323, n41255;
    wire [7:0]\genblk1.write_data_23__N_3541 ;
    wire [7:0]\genblk1.write_data_31__N_3525 ;
    wire [7:0]\genblk1.write_data_15__N_3557 ;
    
    wire n12390;
    wire [31:0]LM32D_DAT_O;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(390[13:24])
    
    wire n41238, n41309, n41461, n10004, n10006, n10008, n41488, 
        n10012, n41485, n10016, n10018, n41482, n10022, n10024, 
        n10026, n10028, n41221, n5_adj_6525, n35788, n15_adj_6526, 
        n41222, n11831, n41307, n41306, n33, n71, n21_adj_6527, 
        LM32D_WE_O, n45079, n45080;
    wire [1:0]selected_1__N_354;
    
    wire LM32D_STB_O, bus_error_f_N_1884, n41429;
    wire [2:0]next_cycle_type;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(347[24:39])
    
    wire n30900, n41410, REF_CLK_c_enable_97;
    wire [31:0]ROM_DAT_O;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(392[26:35])
    wire [31:0]data;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(105[23:27])
    wire [7:0]n69;
    
    wire n33294, n33370, n33256, n33218, n33180, write_enable;
    wire [1:0]state_1__N_3407;
    
    wire n6362;
    wire [7:0]n87;
    
    wire n41289;
    wire [1:0]selected_c;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(244[15:23])
    wire [7:0]n78;
    
    wire n41326, REF_CLK_c_enable_1221;
    wire [3:0]LM32D_SEL_O;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(392[12:23])
    
    wire n41243, REF_CLK_c_enable_1581;
    wire [2:0]LM32I_CTI_O;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(384[12:23])
    
    wire REF_CLK_c_enable_1597, REF_CLK_c_enable_1605, REF_CLK_c_enable_1589, 
        n41387, n9_adj_6532, REF_CLK_c_enable_1558;
    wire [7:0]n96;
    
    wire REF_CLK_c_enable_1574, n32216, n32220, n41226, REF_CLK_c_enable_1131, 
        REF_CLK_c_enable_1550, REF_CLK_c_enable_1566, n37905, n37904, 
        n37906, n37903, LEDGPIO_ACK_O, n5223, n37955, n37956, n37954, 
        n41250;
    wire [31:0]reg_12;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(106[15:21])
    
    wire n2_adj_6536, n40677, n2_adj_6537, n2_adj_6538, n2_adj_6539, 
        n2_adj_6540, n2_adj_6541, n2_adj_6542, n2_adj_6543, n2_adj_6544, 
        n2_adj_6545, n2_adj_6546, n2_adj_6547, n2_adj_6548, n2_adj_6549, 
        n2_adj_6550, n2_adj_6551, n2_adj_6552, n2_adj_6553, PIO_OUT_7__N_3493, 
        write_ack_N_4033, n35736, n32366, n41258;
    
    LUT4 i11_3_lut (.A(ebrEBR_DAT_O[10]), .B(\genblk1.write_data_d [10]), 
         .C(\genblk1.raw_hazard ), .Z(n9)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut.init = 16'hcaca;
    LUT4 i10_3_lut (.A(ebrEBR_DAT_O[9]), .B(\genblk1.write_data_d [9]), 
         .C(\genblk1.raw_hazard ), .Z(n11)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i10_3_lut.init = 16'hcaca;
    LUT4 i31816_2_lut_3_lut_4_lut (.A(n32332), .B(n41210), .C(n41186), 
         .D(\SHAREDBUS_ADR_I[7] ), .Z(n36988)) /* synthesis lut_function=(!(A+!(B (C+!(D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i31816_2_lut_3_lut_4_lut.init = 16'h4044;
    LUT4 i13661_3_lut (.A(ebrEBR_DAT_O[7]), .B(\genblk1.write_data_d [7]), 
         .C(\genblk1.raw_hazard ), .Z(\genblk1.read_data [7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i13661_3_lut.init = 16'hcaca;
    LUT4 i31171_2_lut_3_lut_4_lut (.A(n32332), .B(n41210), .C(n41186), 
         .D(\SHAREDBUS_ADR_I[7] ), .Z(n36343)) /* synthesis lut_function=(A (C+!(D))+!A !(B+!(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i31171_2_lut_3_lut_4_lut.init = 16'hb0bb;
    LUT4 i13693_3_lut (.A(ebrEBR_DAT_O[6]), .B(\genblk1.write_data_d [6]), 
         .C(\genblk1.raw_hazard ), .Z(\genblk1.read_data [6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i13693_3_lut.init = 16'hcaca;
    LUT4 i13102_3_lut (.A(ebrEBR_DAT_O[24]), .B(\genblk1.write_data_d [24]), 
         .C(\genblk1.raw_hazard ), .Z(\genblk1.read_data [24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i13102_3_lut.init = 16'hcaca;
    LUT4 i22488_1_lut (.A(n3), .Z(n1[0])) /* synthesis lut_function=(!(A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(472[15:29])
    defparam i22488_1_lut.init = 16'h5555;
    LUT4 i30706_3_lut_4_lut (.A(n41276), .B(n41253), .C(n32798), .D(n35761), 
         .Z(n35868)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i30706_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_rep_163_2_lut_4_lut (.A(n41234), .B(SHAREDBUS_ADR_I[31]), .C(\SHAREDBUS_ADR_I[10] ), 
         .D(n32332), .Z(n37927)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_rep_163_2_lut_4_lut.init = 16'hfffb;
    LUT4 i1_rep_167_2_lut_4_lut (.A(n41234), .B(SHAREDBUS_ADR_I[31]), .C(\SHAREDBUS_ADR_I[10] ), 
         .D(n32332), .Z(n37931)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_rep_167_2_lut_4_lut.init = 16'hfffb;
    LUT4 i1_rep_166_2_lut_4_lut (.A(n41234), .B(SHAREDBUS_ADR_I[31]), .C(\SHAREDBUS_ADR_I[10] ), 
         .D(n32332), .Z(n37930)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_rep_166_2_lut_4_lut.init = 16'hfffb;
    LUT4 i1_rep_165_2_lut_4_lut (.A(n41234), .B(SHAREDBUS_ADR_I[31]), .C(\SHAREDBUS_ADR_I[10] ), 
         .D(n32332), .Z(n37929)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_rep_165_2_lut_4_lut.init = 16'hfffb;
    LUT4 i1_rep_164_2_lut_4_lut (.A(n41234), .B(SHAREDBUS_ADR_I[31]), .C(\SHAREDBUS_ADR_I[10] ), 
         .D(n32332), .Z(n37928)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_rep_164_2_lut_4_lut.init = 16'hfffb;
    LUT4 i1_2_lut_rep_784_4_lut (.A(n41234), .B(SHAREDBUS_ADR_I[31]), .C(\SHAREDBUS_ADR_I[10] ), 
         .D(n32332), .Z(n41189)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_2_lut_rep_784_4_lut.init = 16'hfffb;
    LUT4 i1_rep_162_2_lut_4_lut (.A(n41234), .B(SHAREDBUS_ADR_I[31]), .C(\SHAREDBUS_ADR_I[10] ), 
         .D(n32332), .Z(n37926)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_rep_162_2_lut_4_lut.init = 16'hfffb;
    LUT4 i1_rep_168_2_lut_4_lut (.A(n41234), .B(SHAREDBUS_ADR_I[31]), .C(\SHAREDBUS_ADR_I[10] ), 
         .D(n32332), .Z(n37932)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_rep_168_2_lut_4_lut.init = 16'hfffb;
    LUT4 i33102_2_lut_4_lut (.A(n41234), .B(SHAREDBUS_ADR_I[31]), .C(\SHAREDBUS_ADR_I[10] ), 
         .D(n41251), .Z(n33368)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i33102_2_lut_4_lut.init = 16'h0004;
    LUT4 i30678_3_lut_4_lut (.A(n41273), .B(n41269), .C(n41277), .D(n41242), 
         .Z(n35840)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30678_3_lut_4_lut.init = 16'hfffe;
    LUT4 i30728_3_lut_4_lut (.A(n41273), .B(n41269), .C(n35712), .D(n15), 
         .Z(n35890)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30728_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut (.A(n41347), .B(n41303), .C(n41246), .D(n41279), 
         .Z(n34698)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0010;
    LUT4 i12_3_lut (.A(n9_adj_6341), .B(\genblk1.EBR_DAT_I_d [19]), .C(\genblk1.EBR_SEL_I_d [2]), 
         .Z(\genblk1.write_data_23__N_3549 [3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i12_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut (.A(n41277), .B(n41236), .C(n33088), .D(n4865[4]), 
         .Z(n32980)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_3_lut_4_lut_adj_746 (.A(n41277), .B(n41236), .C(n33088), .D(n4865[14]), 
         .Z(n32940)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_adj_746.init = 16'h1000;
    LUT4 i1_3_lut_4_lut_adj_747 (.A(n41277), .B(n41236), .C(n33088), .D(n4865[17]), 
         .Z(n33100)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_adj_747.init = 16'h1000;
    LUT4 i1_3_lut_4_lut_adj_748 (.A(n41277), .B(n41236), .C(n33088), .D(n4865[22]), 
         .Z(n33060)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_adj_748.init = 16'h1000;
    LUT4 i1_3_lut_4_lut_adj_749 (.A(n41277), .B(n41236), .C(n33088), .D(n4865[24]), 
         .Z(n32864)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_adj_749.init = 16'h1000;
    FD1P3DX counter_2248__i0 (.D(n1[0]), .SP(REF_CLK_c_enable_1606), .CK(REF_CLK_c), 
            .CD(n41434), .Q(n3));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(472[15:29])
    defparam counter_2248__i0.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut_adj_750 (.A(n41277), .B(n41236), .C(n33088), .D(n4865[29]), 
         .Z(n33020)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_adj_750.init = 16'h1000;
    LUT4 i11_3_lut_adj_751 (.A(n11_adj_6342), .B(\genblk1.EBR_DAT_I_d [21]), 
         .C(\genblk1.EBR_SEL_I_d [2]), .Z(\genblk1.write_data_23__N_3549 [5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_751.init = 16'hcaca;
    LUT4 i12_3_lut_adj_752 (.A(n9_adj_6343), .B(\genblk1.EBR_DAT_I_d [22]), 
         .C(\genblk1.EBR_SEL_I_d [2]), .Z(\genblk1.write_data_23__N_3549 [6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i12_3_lut_adj_752.init = 16'hcaca;
    LUT4 i12_3_lut_adj_753 (.A(n9_adj_6344), .B(\genblk1.EBR_DAT_I_d [23]), 
         .C(\genblk1.EBR_SEL_I_d [2]), .Z(\genblk1.write_data_23__N_3549 [7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i12_3_lut_adj_753.init = 16'hcaca;
    LUT4 i1_4_lut (.A(n34704), .B(n41210), .C(n35633), .D(n34702), .Z(inst1_FIFOof_wr)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_4_lut.init = 16'h0800;
    LUT4 i1_4_lut_adj_754 (.A(n41277), .B(n19), .C(n34692), .D(n41276), 
         .Z(n34704)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_754.init = 16'h0010;
    LUT4 i1_4_lut_adj_755 (.A(n34698), .B(SHAREDBUS_ADR_I[20]), .C(n32798), 
         .D(SHAREDBUS_ADR_I[27]), .Z(n34702)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_755.init = 16'h0002;
    LUT4 i1_4_lut_adj_756 (.A(SHAREDBUS_ADR_I[24]), .B(n41237), .C(n41278), 
         .D(n34672), .Z(n34692)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_756.init = 16'h1000;
    LUT4 i1_3_lut (.A(n41301), .B(n41310), .C(inst3_Full), .Z(n34672)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_3_lut.init = 16'h0808;
    LUT4 i1_4_lut_adj_757 (.A(n31779), .B(n41210), .C(n34664), .D(n35908), 
         .Z(inst1_FIFOif_rd)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_adj_757.init = 16'h0040;
    LUT4 i1_4_lut_adj_758 (.A(n34650), .B(n41225), .C(n19), .D(n35647), 
         .Z(n34664)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_758.init = 16'h0002;
    LUT4 i30746_4_lut (.A(n15), .B(n35796), .C(n41273), .D(n41272), 
         .Z(n35908)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30746_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_759 (.A(n41274), .B(n41246), .C(n34632), .D(n41310), 
         .Z(n34650)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_759.init = 16'h4000;
    LUT4 i1_3_lut_adj_760 (.A(n41301), .B(inst3_Empty), .C(fiford_reg), 
         .Z(n34632)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i1_3_lut_adj_760.init = 16'h0202;
    LUT4 i14544_2_lut_3_lut_4_lut (.A(n41298), .B(SHAREDBUS_ADR_I[15]), 
         .C(n41300), .D(n11769), .Z(n19808)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i14544_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_789_3_lut (.A(n41298), .B(SHAREDBUS_ADR_I[15]), .C(n11769), 
         .Z(n41194)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_2_lut_rep_789_3_lut.init = 16'hfefe;
    LUT4 i33219_3_lut_rep_805_4_lut (.A(n41298), .B(SHAREDBUS_ADR_I[15]), 
         .C(\SHAREDBUS_ADR_I[10] ), .D(SHAREDBUS_ADR_I[31]), .Z(n41210)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i33219_3_lut_rep_805_4_lut.init = 16'h0100;
    LUT4 i1_rep_143_2_lut_3_lut (.A(n41298), .B(SHAREDBUS_ADR_I[15]), .C(n11769), 
         .Z(n37907)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_rep_143_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_rep_145_2_lut_3_lut (.A(n41298), .B(SHAREDBUS_ADR_I[15]), .C(n11769), 
         .Z(n37909)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_rep_145_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_761 (.A(n35942), .B(n31833), .C(SHAREDBUS_ADR_I[31]), 
         .D(n61), .Z(n31955)) /* synthesis lut_function=(!(A+!(B+!(C+!(D))))) */ ;
    defparam i1_4_lut_adj_761.init = 16'h4544;
    LUT4 i30780_4_lut (.A(n35844), .B(n35712), .C(n35888), .D(n41259), 
         .Z(n35942)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30780_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_762 (.A(n35886), .B(n41303), .C(n32728), .D(n41298), 
         .Z(n31833)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_762.init = 16'h0010;
    LUT4 i30726_3_lut (.A(SHAREDBUS_ADR_I[25]), .B(n29), .C(n19), .Z(n35888)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i30726_3_lut.init = 16'hfefe;
    LUT4 i30724_4_lut (.A(n41300), .B(n41301), .C(SHAREDBUS_ADR_I[15]), 
         .D(\SHAREDBUS_ADR_I[10] ), .Z(n35886)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30724_4_lut.init = 16'hfffe;
    LUT4 i33334_4_lut (.A(n32900), .B(n41210), .C(n41262), .D(n32898), 
         .Z(n30762)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i33334_4_lut.init = 16'h0040;
    LUT4 i1_4_lut_adj_763 (.A(n19), .B(n41225), .C(n41263), .D(n32882), 
         .Z(n32900)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_763.init = 16'hfffe;
    LUT4 i1_4_lut_adj_764 (.A(n15), .B(n41265), .C(n32890), .D(n41264), 
         .Z(n32898)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_764.init = 16'hfffe;
    LUT4 i1_2_lut (.A(SHAREDBUS_ADR_I[16]), .B(SHAREDBUS_ADR_I[27]), .Z(n32882)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i33223_4_lut (.A(n32200), .B(n41210), .C(n32194), .D(n19), 
         .Z(REF_CLK_c_enable_424)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i33223_4_lut.init = 16'h0004;
    LUT4 i1_4_lut_adj_765 (.A(n15), .B(n41268), .C(n32192), .D(n41267), 
         .Z(n32200)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_765.init = 16'hfffe;
    LUT4 i1_4_lut_adj_766 (.A(n41269), .B(n41303), .C(n32174), .D(n41301), 
         .Z(n32194)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_766.init = 16'hfffe;
    LUT4 i1_rep_146_2_lut_3_lut (.A(n41298), .B(SHAREDBUS_ADR_I[15]), .C(n11769), 
         .Z(n37910)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_rep_146_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_rep_147_2_lut_3_lut (.A(n41298), .B(SHAREDBUS_ADR_I[15]), .C(n11769), 
         .Z(n37911)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_rep_147_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_rep_144_2_lut_3_lut (.A(n41298), .B(SHAREDBUS_ADR_I[15]), .C(n11769), 
         .Z(n37908)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_rep_144_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_rep_148_2_lut_3_lut (.A(n41298), .B(SHAREDBUS_ADR_I[15]), .C(n11769), 
         .Z(n37912)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_rep_148_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_rep_149_2_lut_3_lut (.A(n41298), .B(SHAREDBUS_ADR_I[15]), .C(n11769), 
         .Z(n37913)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_rep_149_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_830 (.A(SHAREDBUS_ADR_I[16]), .B(SHAREDBUS_ADR_I[20]), 
         .Z(n41235)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_rep_830.init = 16'heeee;
    LUT4 i1_2_lut_3_lut (.A(SHAREDBUS_ADR_I[16]), .B(SHAREDBUS_ADR_I[20]), 
         .C(n41303), .Z(n32028)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_831 (.A(SHAREDBUS_ADR_I[18]), .B(\SHAREDBUS_ADR_I[29] ), 
         .Z(n41236)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_rep_831.init = 16'heeee;
    LUT4 i1_2_lut_rep_832 (.A(SHAREDBUS_ADR_I[30]), .B(SHAREDBUS_ADR_I[25]), 
         .Z(n41237)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_rep_832.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(SHAREDBUS_ADR_I[30]), .B(SHAREDBUS_ADR_I[25]), 
         .C(\SHAREDBUS_ADR_I[29] ), .D(SHAREDBUS_ADR_I[18]), .Z(n32032)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut_adj_767 (.A(SHAREDBUS_ADR_I[30]), .B(SHAREDBUS_ADR_I[25]), 
         .C(n41246), .D(SHAREDBUS_ADR_I[24]), .Z(n35186)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_3_lut_4_lut_adj_767.init = 16'h0010;
    LUT4 i13766_3_lut (.A(ebrEBR_DAT_O[4]), .B(\genblk1.write_data_d [4]), 
         .C(\genblk1.raw_hazard ), .Z(\genblk1.read_data [4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i13766_3_lut.init = 16'hcaca;
    LUT4 i30646_3_lut_4_lut (.A(SHAREDBUS_ADR_I[30]), .B(SHAREDBUS_ADR_I[25]), 
         .C(n41347), .D(\SHAREDBUS_ADR_I[23] ), .Z(n35808)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i30646_3_lut_4_lut.init = 16'hfffe;
    PFUMX i34381 (.BLUT(n41492), .ALUT(n41493), .C0(n45101), .Z(n19));
    LUT4 i1_4_lut_adj_768 (.A(n41220), .B(n32694), .C(n19), .D(n32690), 
         .Z(n11769)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_768.init = 16'hfffe;
    LUT4 i1_4_lut_rep_788 (.A(n35912), .B(n41210), .C(n35633), .D(n32464), 
         .Z(n41193)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_rep_788.init = 16'h0400;
    LUT4 i1_4_lut_adj_769 (.A(n41274), .B(n29), .C(SHAREDBUS_ADR_I[18]), 
         .D(SHAREDBUS_ADR_I[31]), .Z(n32694)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_769.init = 16'hfffe;
    LUT4 i1_2_lut_rep_790 (.A(SHAREDBUS_ADR_I[15]), .B(n11769), .Z(n41195)) /* synthesis lut_function=((B)+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_rep_790.init = 16'hdddd;
    LUT4 mux_65_i1_3_lut_3_lut_4_lut (.A(SHAREDBUS_ADR_I[15]), .B(n11769), 
         .C(n1030[0]), .D(ebrEBR_ACK_O), .Z(n1063[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam mux_65_i1_3_lut_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i31_3_lut_3_lut_4_lut (.A(SHAREDBUS_ADR_I[15]), .B(n11769), .C(n21), 
         .D(ebrEBR_DAT_O[24]), .Z(n16)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i31_3_lut_3_lut_4_lut.init = 16'hf2d0;
    FD1S3DX counter_2248__i2 (.D(n12428), .CK(REF_CLK_c), .CD(n41434), 
            .Q(\counter[2] ));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(472[15:29])
    defparam counter_2248__i2.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_770 (.A(n34992), .B(REF_CLK_c_enable_424), .C(n41310), 
         .D(n41346), .Z(PIO_DATAI_0__N_3822)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_770.init = 16'h0008;
    FD1P3DX counter_2248__i1 (.D(n1[1]), .SP(REF_CLK_c_enable_1606), .CK(REF_CLK_c), 
            .CD(n41434), .Q(n2));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(472[15:29])
    defparam counter_2248__i1.GSR = "ENABLED";
    LUT4 i11_3_lut_adj_771 (.A(n11), .B(\genblk1.EBR_DAT_I_d [9]), .C(\genblk1.EBR_SEL_I_d [1]), 
         .Z(\genblk1.write_data_15__N_3565 [1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_771.init = 16'hcaca;
    LUT4 i12_3_lut_adj_772 (.A(n9), .B(\genblk1.EBR_DAT_I_d [10]), .C(\genblk1.EBR_SEL_I_d [1]), 
         .Z(\genblk1.write_data_15__N_3565 [2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i12_3_lut_adj_772.init = 16'hcaca;
    LUT4 i11_3_lut_adj_773 (.A(n11_adj_6346), .B(\genblk1.EBR_DAT_I_d [11]), 
         .C(\genblk1.EBR_SEL_I_d [1]), .Z(\genblk1.write_data_15__N_3565 [3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_773.init = 16'hcaca;
    LUT4 i13801_3_lut (.A(ebrEBR_DAT_O[3]), .B(\genblk1.write_data_d [3]), 
         .C(\genblk1.raw_hazard ), .Z(\genblk1.read_data [3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i13801_3_lut.init = 16'hcaca;
    LUT4 mux_67_i1_4_lut (.A(spiSPI_ACK_O), .B(n32084), .C(n47), .D(n41210), 
         .Z(n997[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(554[1] 556[2])
    defparam mux_67_i1_4_lut.init = 16'hca0a;
    LUT4 i32946_4_lut (.A(n997[0]), .B(n1096[0]), .C(n41194), .D(n41181), 
         .Z(SHAREDBUS_ACK_O_N_91[0])) /* synthesis lut_function=(A (B+(C (D)))+!A !((C (D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(549[1] 556[2])
    defparam i32946_4_lut.init = 16'haccc;
    LUT4 i13617_4_lut (.A(spiSPI_DAT_O[9]), .B(FIFOwb_en), .C(n47), .D(FIFOwb_DAT_O[9]), 
         .Z(n3_adj_6347)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i13617_4_lut.init = 16'hca0a;
    LUT4 i13_4_lut (.A(n34304), .B(reg_00[9]), .C(n41185), .D(n34226), 
         .Z(n15_adj_6348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i13_4_lut.init = 16'hcfca;
    LUT4 i13547_4_lut (.A(spiSPI_DAT_O[11]), .B(FIFOwb_en), .C(n47), .D(FIFOwb_DAT_O[11]), 
         .Z(n3_adj_6349)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i13547_4_lut.init = 16'hca0a;
    LUT4 i13_4_lut_adj_774 (.A(n34304), .B(reg_00[11]), .C(n41185), .D(n34302), 
         .Z(n15_adj_6350)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i13_4_lut_adj_774.init = 16'hcfca;
    LUT4 i13477_4_lut (.A(spiSPI_DAT_O[13]), .B(FIFOwb_en), .C(n47), .D(FIFOwb_DAT_O[13]), 
         .Z(n3_adj_6351)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i13477_4_lut.init = 16'hca0a;
    LUT4 i13_4_lut_adj_775 (.A(n34304), .B(reg_00[13]), .C(n41185), .D(n34378), 
         .Z(n15_adj_6352)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i13_4_lut_adj_775.init = 16'hcfca;
    LUT4 i13407_4_lut (.A(spiSPI_DAT_O[15]), .B(FIFOwb_en), .C(n47), .D(FIFOwb_DAT_O[15]), 
         .Z(n3_adj_6353)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i13407_4_lut.init = 16'hca0a;
    LUT4 i13_4_lut_adj_776 (.A(n34304), .B(reg_00[15]), .C(n41185), .D(n34416), 
         .Z(n15_adj_6354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i13_4_lut_adj_776.init = 16'hcfca;
    LUT4 i12_3_lut_adj_777 (.A(n9_adj_6355), .B(\genblk1.EBR_DAT_I_d [12]), 
         .C(\genblk1.EBR_SEL_I_d [1]), .Z(\genblk1.write_data_15__N_3565 [4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i12_3_lut_adj_777.init = 16'hcaca;
    LUT4 i12949_4_lut (.A(spiSPI_DAT_O[28]), .B(FIFOwb_en), .C(n47), .D(FIFOwb_DAT_O[28]), 
         .Z(n3_adj_6356)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i12949_4_lut.init = 16'hca0a;
    LUT4 i13_4_lut_adj_778 (.A(n34304), .B(reg_00[28]), .C(n41185), .D(n34340), 
         .Z(n15_adj_6357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i13_4_lut_adj_778.init = 16'hcfca;
    LUT4 i13196_4_lut (.A(spiSPI_DAT_O[21]), .B(FIFOwb_en), .C(n47), .D(FIFOwb_DAT_O[21]), 
         .Z(n3_adj_6358)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i13196_4_lut.init = 16'hca0a;
    LUT4 i13_4_lut_adj_779 (.A(n34304), .B(reg_00[21]), .C(n41185), .D(n34264), 
         .Z(n15_adj_6359)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i13_4_lut_adj_779.init = 16'hcfca;
    LUT4 i7_4_lut (.A(spiSPI_DAT_O[29]), .B(n33030), .C(n47), .D(n30762), 
         .Z(n17)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'hca0a;
    LUT4 i12910_4_lut (.A(n33368), .B(reg_00[29]), .C(n41185), .D(n33366), 
         .Z(n13)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i12910_4_lut.init = 16'hcac0;
    LUT4 i13055_4_lut (.A(spiSPI_DAT_O[25]), .B(FIFOwb_en), .C(n47), .D(FIFOwb_DAT_O[25]), 
         .Z(n3_adj_6360)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i13055_4_lut.init = 16'hca0a;
    LUT4 i13_4_lut_adj_780 (.A(n34304), .B(reg_00[25]), .C(n41185), .D(n34036), 
         .Z(n15_adj_6361)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i13_4_lut_adj_780.init = 16'hcfca;
    LUT4 i13301_4_lut (.A(spiSPI_DAT_O[18]), .B(FIFOwb_en), .C(n47), .D(FIFOwb_DAT_O[18]), 
         .Z(n3_adj_6362)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i13301_4_lut.init = 16'hca0a;
    LUT4 i13_4_lut_adj_781 (.A(n34304), .B(reg_00[18]), .C(n41185), .D(n34188), 
         .Z(n15_adj_6363)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i13_4_lut_adj_781.init = 16'hcfca;
    LUT4 i17_4_lut (.A(spiSPI_DAT_O[24]), .B(n32874), .C(n47), .D(n30762), 
         .Z(n23)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i17_4_lut.init = 16'hca0a;
    LUT4 i7_4_lut_adj_782 (.A(spiSPI_DAT_O[22]), .B(n33070), .C(n47), 
         .D(n30762), .Z(n17_adj_6364)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_782.init = 16'hca0a;
    LUT4 i13157_4_lut (.A(n33368), .B(reg_00[22]), .C(n41185), .D(n33252), 
         .Z(n13_adj_6365)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i13157_4_lut.init = 16'hcac0;
    LUT4 i7_4_lut_adj_783 (.A(spiSPI_DAT_O[17]), .B(n33110), .C(n47), 
         .D(n30762), .Z(n17_adj_6366)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_783.init = 16'hca0a;
    LUT4 i13332_4_lut (.A(n33368), .B(reg_00[17]), .C(n41185), .D(n33290), 
         .Z(n13_adj_6367)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i13332_4_lut.init = 16'hcac0;
    LUT4 i7_4_lut_adj_784 (.A(spiSPI_DAT_O[14]), .B(n32950), .C(n47), 
         .D(n30762), .Z(n17_adj_6368)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_784.init = 16'hca0a;
    LUT4 i13438_4_lut (.A(n33368), .B(reg_00[14]), .C(n41185), .D(n33404), 
         .Z(n13_adj_6369)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i13438_4_lut.init = 16'hcac0;
    LUT4 i13654_4_lut (.A(spiSPI_DAT_O[7]), .B(FIFOwb_en), .C(n47), .D(n30944), 
         .Z(n6)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i13654_4_lut.init = 16'hca0a;
    LUT4 i13646_4_lut (.A(n34304), .B(GPOout_pins[7]), .C(n41185), .D(n34150), 
         .Z(n4)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i13646_4_lut.init = 16'hcfca;
    LUT4 i13686_4_lut (.A(spiSPI_DAT_O[6]), .B(FIFOwb_en), .C(n47), .D(n30948), 
         .Z(n6_adj_6370)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i13686_4_lut.init = 16'hca0a;
    LUT4 i13678_4_lut (.A(n34304), .B(GPOout_pins[6]), .C(n41185), .D(n34454), 
         .Z(n4_adj_6371)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i13678_4_lut.init = 16'hcfca;
    LUT4 i7_4_lut_adj_785 (.A(spiSPI_DAT_O[4]), .B(n32990), .C(n47), .D(n30762), 
         .Z(n15_adj_6372)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_785.init = 16'hca0a;
    LUT4 i13751_4_lut (.A(n33368), .B(GPOout_pins[4]), .C(n41185), .D(n33328), 
         .Z(n11_adj_6373)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i13751_4_lut.init = 16'hcac0;
    LUT4 i13794_4_lut (.A(spiSPI_DAT_O[3]), .B(FIFOwb_en), .C(n47), .D(n30951), 
         .Z(n6_adj_6374)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i13794_4_lut.init = 16'hca0a;
    LUT4 i13786_4_lut (.A(n34304), .B(GPOout_pins[3]), .C(n41185), .D(n34074), 
         .Z(n4_adj_6375)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i13786_4_lut.init = 16'hcfca;
    LUT4 i13826_4_lut (.A(spiSPI_DAT_O[2]), .B(FIFOwb_en), .C(n47), .D(n30949), 
         .Z(n6_adj_6376)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i13826_4_lut.init = 16'hca0a;
    LUT4 i13818_4_lut (.A(n34304), .B(GPOout_pins[2]), .C(n41185), .D(n33998), 
         .Z(n4_adj_6377)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i13818_4_lut.init = 16'hcfca;
    LUT4 mux_107_i1_4_lut (.A(spiSPI_DAT_O[0]), .B(FIFOwb_DAT_O[0]), .C(n47), 
         .D(FIFOwb_en), .Z(n295[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(536[1] 538[2])
    defparam mux_107_i1_4_lut.init = 16'hca0a;
    LUT4 mux_107_i2_4_lut (.A(spiSPI_DAT_O[1]), .B(FIFOwb_DAT_O[1]), .C(n47), 
         .D(FIFOwb_en), .Z(n295[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(536[1] 538[2])
    defparam mux_107_i2_4_lut.init = 16'hca0a;
    LUT4 mux_107_i6_4_lut (.A(spiSPI_DAT_O[5]), .B(FIFOwb_DAT_O[5]), .C(n47), 
         .D(FIFOwb_en), .Z(n295[5])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(536[1] 538[2])
    defparam mux_107_i6_4_lut.init = 16'hca0a;
    LUT4 mux_107_i9_4_lut (.A(spiSPI_DAT_O[8]), .B(FIFOwb_DAT_O[8]), .C(n47), 
         .D(FIFOwb_en), .Z(n295[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(536[1] 538[2])
    defparam mux_107_i9_4_lut.init = 16'hca0a;
    LUT4 i11_3_lut_adj_786 (.A(n11_adj_6378), .B(\genblk1.EBR_DAT_I_d [13]), 
         .C(\genblk1.EBR_SEL_I_d [1]), .Z(\genblk1.write_data_15__N_3565 [5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_786.init = 16'hcaca;
    LUT4 i6_4_lut (.A(spiSPI_DAT_O[31]), .B(FIFOwb_en), .C(n47), .D(FIFOwb_DAT_O[31]), 
         .Z(n17_adj_6379)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'hca0a;
    LUT4 i7_4_lut_adj_787 (.A(spiSPI_DAT_O[30]), .B(FIFOwb_en), .C(n47), 
         .D(FIFOwb_DAT_O[30]), .Z(n17_adj_6380)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_787.init = 16'hca0a;
    LUT4 i7_4_lut_adj_788 (.A(spiSPI_DAT_O[27]), .B(FIFOwb_en), .C(n47), 
         .D(FIFOwb_DAT_O[27]), .Z(n17_adj_6381)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_788.init = 16'hca0a;
    LUT4 i7_4_lut_adj_789 (.A(spiSPI_DAT_O[26]), .B(FIFOwb_en), .C(n47), 
         .D(FIFOwb_DAT_O[26]), .Z(n17_adj_6382)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_789.init = 16'hca0a;
    LUT4 i7_4_lut_adj_790 (.A(spiSPI_DAT_O[23]), .B(FIFOwb_en), .C(n47), 
         .D(FIFOwb_DAT_O[23]), .Z(n17_adj_6383)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_790.init = 16'hca0a;
    LUT4 i7_4_lut_adj_791 (.A(spiSPI_DAT_O[20]), .B(FIFOwb_DAT_O[20]), .C(n47), 
         .D(FIFOwb_en), .Z(n15_adj_6384)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_791.init = 16'hca0a;
    LUT4 i7_4_lut_adj_792 (.A(spiSPI_DAT_O[19]), .B(FIFOwb_en), .C(n47), 
         .D(FIFOwb_DAT_O[19]), .Z(n17_adj_6385)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_792.init = 16'hca0a;
    LUT4 i7_4_lut_adj_793 (.A(spiSPI_DAT_O[16]), .B(FIFOwb_en), .C(n47), 
         .D(FIFOwb_DAT_O[16]), .Z(n17_adj_6386)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_793.init = 16'hca0a;
    LUT4 i7_4_lut_adj_794 (.A(spiSPI_DAT_O[12]), .B(FIFOwb_en), .C(n47), 
         .D(FIFOwb_DAT_O[12]), .Z(n17_adj_6387)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_794.init = 16'hca0a;
    LUT4 i7_4_lut_adj_795 (.A(spiSPI_DAT_O[10]), .B(FIFOwb_en), .C(n47), 
         .D(FIFOwb_DAT_O[10]), .Z(n17_adj_6388)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i7_4_lut_adj_795.init = 16'hca0a;
    LUT4 i1_4_lut_adj_796 (.A(n41181), .B(ebrEBR_DAT_O[9]), .C(n17_adj_6389), 
         .D(n41195), .Z(n14)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_796.init = 16'ha088;
    LUT4 i1_4_lut_adj_797 (.A(n41181), .B(ebrEBR_DAT_O[11]), .C(n17_adj_6390), 
         .D(n41195), .Z(n14_adj_6391)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_797.init = 16'ha088;
    LUT4 i1_4_lut_adj_798 (.A(n41181), .B(ebrEBR_DAT_O[29]), .C(n26), 
         .D(n41195), .Z(n11_adj_6392)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_798.init = 16'ha088;
    LUT4 i1_4_lut_adj_799 (.A(n41181), .B(ebrEBR_DAT_O[13]), .C(n17_adj_6393), 
         .D(n41195), .Z(n14_adj_6394)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_799.init = 16'ha088;
    LUT4 i12_3_lut_adj_800 (.A(n9_adj_6395), .B(\genblk1.EBR_DAT_I_d [14]), 
         .C(\genblk1.EBR_SEL_I_d [1]), .Z(\genblk1.write_data_15__N_3565 [6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i12_3_lut_adj_800.init = 16'hcaca;
    LUT4 i1_4_lut_adj_801 (.A(n41181), .B(ebrEBR_DAT_O[14]), .C(n5), .D(n41195), 
         .Z(n11_adj_6396)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_801.init = 16'ha088;
    LUT4 i1_4_lut_adj_802 (.A(n41181), .B(ebrEBR_DAT_O[15]), .C(n17_adj_6397), 
         .D(n41195), .Z(n14_adj_6398)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_802.init = 16'ha088;
    LUT4 i11_3_lut_adj_803 (.A(n11_adj_6399), .B(\genblk1.EBR_DAT_I_d [15]), 
         .C(\genblk1.EBR_SEL_I_d [1]), .Z(\genblk1.write_data_15__N_3565 [7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_803.init = 16'hcaca;
    LUT4 i11_3_lut_adj_804 (.A(n11_adj_6400), .B(\genblk1.EBR_DAT_I_d [25]), 
         .C(\genblk1.EBR_SEL_I_d [3]), .Z(\genblk1.write_data_31__N_3533 [1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_804.init = 16'hcaca;
    LUT4 i1_4_lut_adj_805 (.A(n949[0]), .B(n30241), .C(n31750), .D(n31955), 
         .Z(n13990)) /* synthesis lut_function=(A+!((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(549[1] 556[2])
    defparam i1_4_lut_adj_805.init = 16'haaae;
    LUT4 i33429_then_3_lut (.A(LM32D_ADR_O[21]), .B(selected[0]), .C(LM32D_ADR_O[28]), 
         .Z(n41493)) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;
    defparam i33429_then_3_lut.init = 16'h3232;
    LUT4 i1_4_lut_adj_806 (.A(n41181), .B(ebrEBR_DAT_O[17]), .C(n5_adj_6401), 
         .D(n41195), .Z(n11_adj_6402)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_806.init = 16'ha088;
    LUT4 i12_3_lut_adj_807 (.A(n9_adj_6403), .B(\genblk1.EBR_DAT_I_d [26]), 
         .C(\genblk1.EBR_SEL_I_d [3]), .Z(\genblk1.write_data_31__N_3533 [2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i12_3_lut_adj_807.init = 16'hcaca;
    LUT4 i1_4_lut_adj_808 (.A(n41181), .B(ebrEBR_DAT_O[18]), .C(n22), 
         .D(n41195), .Z(n9_adj_6404)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_808.init = 16'ha088;
    LUT4 i1_4_lut_adj_809 (.A(n41181), .B(ebrEBR_DAT_O[25]), .C(n22_adj_6405), 
         .D(n41195), .Z(n9_adj_6406)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_809.init = 16'ha088;
    LUT4 i33429_else_3_lut (.A(LM32I_ADR_O[28]), .B(LM32I_ADR_O[21]), .C(selected[0]), 
         .Z(n41492)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i33429_else_3_lut.init = 16'he0e0;
    LUT4 i1_4_lut_adj_810 (.A(n41181), .B(ebrEBR_DAT_O[21]), .C(n22_adj_6407), 
         .D(n41195), .Z(n9_adj_6408)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_810.init = 16'ha088;
    LUT4 i1_4_lut_adj_811 (.A(n41181), .B(ebrEBR_DAT_O[2]), .C(n2_adj_6409), 
         .D(n41195), .Z(n11_adj_6410)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_811.init = 16'ha088;
    LUT4 i1_4_lut_adj_812 (.A(n41181), .B(ebrEBR_DAT_O[3]), .C(n2_adj_6411), 
         .D(n41195), .Z(n11_adj_6412)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_812.init = 16'ha088;
    LUT4 i1_4_lut_adj_813 (.A(n41181), .B(ebrEBR_DAT_O[28]), .C(n22_adj_6413), 
         .D(n41195), .Z(n9_adj_6414)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_813.init = 16'ha088;
    LUT4 i1_4_lut_adj_814 (.A(n41181), .B(ebrEBR_DAT_O[4]), .C(n5_adj_6415), 
         .D(n41195), .Z(n11_adj_6416)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_814.init = 16'ha088;
    LUT4 i1_4_lut_adj_815 (.A(n41181), .B(ebrEBR_DAT_O[6]), .C(n2_adj_6417), 
         .D(n41195), .Z(n11_adj_6418)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_815.init = 16'ha088;
    LUT4 i1_4_lut_adj_816 (.A(n41181), .B(ebrEBR_DAT_O[22]), .C(n26_adj_6419), 
         .D(n41195), .Z(n11_adj_6420)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_816.init = 16'ha088;
    LUT4 i1_4_lut_adj_817 (.A(n41181), .B(ebrEBR_DAT_O[7]), .C(n2_adj_6421), 
         .D(n41195), .Z(n11_adj_6422)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_817.init = 16'ha088;
    LUT4 i1_4_lut_adj_818 (.A(n41181), .B(ebrEBR_DAT_O[0]), .C(n361[0]), 
         .D(n41195), .Z(n11_adj_6423)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(531[1] 538[2])
    defparam i1_4_lut_adj_818.init = 16'ha088;
    LUT4 i1_4_lut_adj_819 (.A(n41181), .B(ebrEBR_DAT_O[10]), .C(n5_adj_6424), 
         .D(n41195), .Z(n11_adj_6425)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_819.init = 16'ha088;
    LUT4 i1_4_lut_adj_820 (.A(n41181), .B(ebrEBR_DAT_O[1]), .C(n361[1]), 
         .D(n41195), .Z(n11_adj_6426)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(531[1] 538[2])
    defparam i1_4_lut_adj_820.init = 16'ha088;
    LUT4 i1_4_lut_adj_821 (.A(n41181), .B(ebrEBR_DAT_O[23]), .C(n25), 
         .D(n41195), .Z(n11_adj_6427)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_821.init = 16'ha088;
    LUT4 i1_4_lut_adj_822 (.A(n41181), .B(ebrEBR_DAT_O[12]), .C(n5_adj_6428), 
         .D(n41195), .Z(n11_adj_6429)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_822.init = 16'ha088;
    LUT4 i1_4_lut_adj_823 (.A(n41181), .B(ebrEBR_DAT_O[5]), .C(n361[5]), 
         .D(n41195), .Z(n11_adj_6430)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(531[1] 538[2])
    defparam i1_4_lut_adj_823.init = 16'ha088;
    LUT4 i1_4_lut_adj_824 (.A(n41181), .B(ebrEBR_DAT_O[30]), .C(n25_adj_6431), 
         .D(n41195), .Z(n11_adj_6432)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_824.init = 16'ha088;
    LUT4 i1_4_lut_adj_825 (.A(n41181), .B(ebrEBR_DAT_O[31]), .C(n25_adj_6433), 
         .D(n41195), .Z(n11_adj_6434)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_825.init = 16'ha088;
    LUT4 i1_4_lut_adj_826 (.A(n41181), .B(ebrEBR_DAT_O[16]), .C(n5_adj_6435), 
         .D(n41195), .Z(n11_adj_6436)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_826.init = 16'ha088;
    LUT4 i1_4_lut_adj_827 (.A(n41181), .B(ebrEBR_DAT_O[26]), .C(n25_adj_6437), 
         .D(n41195), .Z(n11_adj_6438)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_827.init = 16'ha088;
    LUT4 i1_4_lut_adj_828 (.A(n41181), .B(ebrEBR_DAT_O[19]), .C(n25_adj_6439), 
         .D(n41195), .Z(n11_adj_6440)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_828.init = 16'ha088;
    LUT4 i1_4_lut_adj_829 (.A(n41181), .B(ebrEBR_DAT_O[20]), .C(n22_adj_6441), 
         .D(n41195), .Z(n11_adj_6442)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_829.init = 16'ha088;
    LUT4 i1_4_lut_adj_830 (.A(n15), .B(n41210), .C(n32038), .D(n32036), 
         .Z(n30986)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_830.init = 16'hfffb;
    LUT4 i1_4_lut_adj_831 (.A(n41181), .B(ebrEBR_DAT_O[27]), .C(n25_adj_6443), 
         .D(n41195), .Z(n11_adj_6444)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_831.init = 16'ha088;
    LUT4 i12_3_lut_adj_832 (.A(n9_adj_6445), .B(\genblk1.EBR_DAT_I_d [27]), 
         .C(\genblk1.EBR_SEL_I_d [3]), .Z(\genblk1.write_data_31__N_3533 [3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i12_3_lut_adj_832.init = 16'hcaca;
    LUT4 i1_4_lut_adj_833 (.A(n41181), .B(ebrEBR_DAT_O[8]), .C(n361[8]), 
         .D(n41195), .Z(n11_adj_6446)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(531[1] 538[2])
    defparam i1_4_lut_adj_833.init = 16'ha088;
    LUT4 i1_4_lut_adj_834 (.A(n35200), .B(n41210), .C(n15), .D(n35892), 
         .Z(n31476)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_834.init = 16'h0008;
    LUT4 i1_4_lut_adj_835 (.A(n35186), .B(n41225), .C(n19), .D(n35184), 
         .Z(n35200)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_835.init = 16'h0200;
    LUT4 i30730_4_lut (.A(n41270), .B(n41266), .C(n41254), .D(n41268), 
         .Z(n35892)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30730_4_lut.init = 16'hfffe;
    LUT4 i11_3_lut_adj_836 (.A(n11_adj_6447), .B(\genblk1.EBR_DAT_I_d [28]), 
         .C(\genblk1.EBR_SEL_I_d [3]), .Z(\genblk1.write_data_31__N_3533 [4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_836.init = 16'hcaca;
    LUT4 i13833_3_lut (.A(ebrEBR_DAT_O[2]), .B(\genblk1.write_data_d [2]), 
         .C(\genblk1.raw_hazard ), .Z(\genblk1.read_data [2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i13833_3_lut.init = 16'hcaca;
    LUT4 i12_3_lut_adj_837 (.A(n9_adj_6448), .B(\genblk1.EBR_DAT_I_d [29]), 
         .C(\genblk1.EBR_SEL_I_d [3]), .Z(\genblk1.write_data_31__N_3533 [5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i12_3_lut_adj_837.init = 16'hcaca;
    LUT4 i12_3_lut_adj_838 (.A(n9_adj_6449), .B(\genblk1.EBR_DAT_I_d [30]), 
         .C(\genblk1.EBR_SEL_I_d [3]), .Z(\genblk1.write_data_31__N_3533 [6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i12_3_lut_adj_838.init = 16'hcaca;
    LUT4 i11_3_lut_adj_839 (.A(n7), .B(\genblk1.EBR_DAT_I_d [31]), .C(\genblk1.EBR_SEL_I_d [3]), 
         .Z(\genblk1.write_data_31__N_3533 [7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_839.init = 16'hcaca;
    LUT4 i12_3_lut_adj_840 (.A(n9_adj_6450), .B(\genblk1.EBR_DAT_I_d [17]), 
         .C(\genblk1.EBR_SEL_I_d [2]), .Z(\genblk1.write_data_23__N_3549 [1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i12_3_lut_adj_840.init = 16'hcaca;
    LUT4 i11_3_lut_adj_841 (.A(n11_adj_6451), .B(\genblk1.EBR_DAT_I_d [18]), 
         .C(\genblk1.EBR_SEL_I_d [2]), .Z(\genblk1.write_data_23__N_3549 [2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_841.init = 16'hcaca;
    LUT4 i11_3_lut_adj_842 (.A(ebrEBR_DAT_O[16]), .B(\genblk1.write_data_d [16]), 
         .C(\genblk1.raw_hazard ), .Z(n9_adj_6452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_842.init = 16'hcaca;
    LUT4 i30750_4_lut (.A(n35796), .B(n19), .C(n35605), .D(n41269), 
         .Z(n35912)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30750_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_843 (.A(n41279), .B(n41236), .C(n33088), .D(n35649), 
         .Z(n32464)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_843.init = 16'h0010;
    LUT4 i30491_2_lut (.A(SHAREDBUS_ADR_I[27]), .B(SHAREDBUS_ADR_I[24]), 
         .Z(n35649)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i30491_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_844 (.A(n35160), .B(n41210), .C(n35890), .D(n41225), 
         .Z(write_ack_N_4649)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_844.init = 16'h0008;
    LUT4 i1_4_lut_adj_845 (.A(n41260), .B(n19), .C(n32312), .D(n35136), 
         .Z(n35160)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_845.init = 16'h0100;
    LUT4 i1_4_lut_adj_846 (.A(n31779), .B(n41210), .C(n35236), .D(n35890), 
         .Z(fiford)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_adj_846.init = 16'h0040;
    LUT4 i1_4_lut_adj_847 (.A(n35222), .B(n41225), .C(n19), .D(n32312), 
         .Z(n35236)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_847.init = 16'h0002;
    LUT4 i1_4_lut_adj_848 (.A(n41260), .B(n41246), .C(n35204), .D(n41310), 
         .Z(n35222)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_848.init = 16'h4000;
    LUT4 i22490_2_lut (.A(n2), .B(n3), .Z(n1[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(472[15:29])
    defparam i22490_2_lut.init = 16'h6666;
    LUT4 i11_3_lut_adj_849 (.A(ebrEBR_DAT_O[23]), .B(\genblk1.write_data_d [23]), 
         .C(\genblk1.raw_hazard ), .Z(n9_adj_6344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_849.init = 16'hcaca;
    LUT4 i11_3_lut_adj_850 (.A(ebrEBR_DAT_O[22]), .B(\genblk1.write_data_d [22]), 
         .C(\genblk1.raw_hazard ), .Z(n9_adj_6343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_850.init = 16'hcaca;
    LUT4 i10_3_lut_adj_851 (.A(ebrEBR_DAT_O[21]), .B(\genblk1.write_data_d [21]), 
         .C(\genblk1.raw_hazard ), .Z(n11_adj_6342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i10_3_lut_adj_851.init = 16'hcaca;
    LUT4 i13241_3_lut (.A(ebrEBR_DAT_O[20]), .B(\genblk1.write_data_d [20]), 
         .C(\genblk1.raw_hazard ), .Z(\genblk1.read_data [20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i13241_3_lut.init = 16'hcaca;
    LUT4 i11_3_lut_adj_852 (.A(ebrEBR_DAT_O[19]), .B(\genblk1.write_data_d [19]), 
         .C(\genblk1.raw_hazard ), .Z(n9_adj_6341)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_852.init = 16'hcaca;
    LUT4 i10_3_lut_adj_853 (.A(ebrEBR_DAT_O[18]), .B(\genblk1.write_data_d [18]), 
         .C(\genblk1.raw_hazard ), .Z(n11_adj_6451)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i10_3_lut_adj_853.init = 16'hcaca;
    LUT4 i11_3_lut_adj_854 (.A(ebrEBR_DAT_O[17]), .B(\genblk1.write_data_d [17]), 
         .C(\genblk1.raw_hazard ), .Z(n9_adj_6450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_854.init = 16'hcaca;
    LUT4 i10_3_lut_adj_855 (.A(ebrEBR_DAT_O[31]), .B(\genblk1.write_data_d [31]), 
         .C(\genblk1.raw_hazard ), .Z(n7)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i10_3_lut_adj_855.init = 16'hcaca;
    LUT4 i11_3_lut_adj_856 (.A(ebrEBR_DAT_O[30]), .B(\genblk1.write_data_d [30]), 
         .C(\genblk1.raw_hazard ), .Z(n9_adj_6449)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_856.init = 16'hcaca;
    LUT4 i11_3_lut_adj_857 (.A(ebrEBR_DAT_O[29]), .B(\genblk1.write_data_d [29]), 
         .C(\genblk1.raw_hazard ), .Z(n9_adj_6448)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_857.init = 16'hcaca;
    LUT4 i10_3_lut_adj_858 (.A(ebrEBR_DAT_O[28]), .B(\genblk1.write_data_d [28]), 
         .C(\genblk1.raw_hazard ), .Z(n11_adj_6447)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i10_3_lut_adj_858.init = 16'hcaca;
    LUT4 i11_3_lut_adj_859 (.A(ebrEBR_DAT_O[27]), .B(\genblk1.write_data_d [27]), 
         .C(\genblk1.raw_hazard ), .Z(n9_adj_6445)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_859.init = 16'hcaca;
    LUT4 i11_3_lut_adj_860 (.A(ebrEBR_DAT_O[26]), .B(\genblk1.write_data_d [26]), 
         .C(\genblk1.raw_hazard ), .Z(n9_adj_6403)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_860.init = 16'hcaca;
    LUT4 i10_3_lut_adj_861 (.A(ebrEBR_DAT_O[25]), .B(\genblk1.write_data_d [25]), 
         .C(\genblk1.raw_hazard ), .Z(n11_adj_6400)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i10_3_lut_adj_861.init = 16'hcaca;
    LUT4 i10_3_lut_adj_862 (.A(ebrEBR_DAT_O[15]), .B(\genblk1.write_data_d [15]), 
         .C(\genblk1.raw_hazard ), .Z(n11_adj_6399)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i10_3_lut_adj_862.init = 16'hcaca;
    LUT4 i1_3_lut_rep_847 (.A(n954[0]), .B(\SHAREDBUS_ADR_I[7] ), .C(GPIOGPIO_ACK_O), 
         .Z(n41252)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_3_lut_rep_847.init = 16'h0808;
    LUT4 i1_4_lut_adj_863 (.A(\SHAREDBUS_ADR_I[5] ), .B(n41310), .C(n41346), 
         .D(n34960), .Z(n34966)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_863.init = 16'h0100;
    LUT4 i1_3_lut_adj_864 (.A(n954[0]), .B(\SHAREDBUS_ADR_I[7] ), .C(GPIOGPIO_ACK_O), 
         .Z(n34960)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_864.init = 16'h8080;
    LUT4 i11_3_lut_adj_865 (.A(ebrEBR_DAT_O[14]), .B(\genblk1.write_data_d [14]), 
         .C(\genblk1.raw_hazard ), .Z(n9_adj_6395)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_865.init = 16'hcaca;
    LUT4 i1_4_lut_adj_866 (.A(n41275), .B(n41310), .C(n41239), .D(n41252), 
         .Z(n34926)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_866.init = 16'h1000;
    LUT4 i1_2_lut_4_lut_adj_867 (.A(n954[0]), .B(\SHAREDBUS_ADR_I[7] ), 
         .C(GPIOGPIO_ACK_O), .D(\SHAREDBUS_ADR_I[5] ), .Z(n34992)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_867.init = 16'h0008;
    LUT4 i10_3_lut_adj_868 (.A(ebrEBR_DAT_O[13]), .B(\genblk1.write_data_d [13]), 
         .C(\genblk1.raw_hazard ), .Z(n11_adj_6378)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i10_3_lut_adj_868.init = 16'hcaca;
    LUT4 i1_2_lut_rep_848 (.A(SHAREDBUS_ADR_I[20]), .B(\SHAREDBUS_ADR_I[22] ), 
         .Z(n41253)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_rep_848.init = 16'heeee;
    LUT4 i32986_4_lut (.A(n31), .B(n16), .C(n41195), .D(n36988), .Z(n13_adj_6453)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;
    defparam i32986_4_lut.init = 16'hccac;
    LUT4 i1_4_lut_adj_869 (.A(n32326), .B(n34372), .C(n32322), .D(n19), 
         .Z(n32332)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_869.init = 16'hfffe;
    LUT4 i1_4_lut_adj_870 (.A(n15), .B(n32304), .C(n32312), .D(n41310), 
         .Z(n32326)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_870.init = 16'hfffe;
    LUT4 i1_4_lut_adj_871 (.A(n32318), .B(SHAREDBUS_ADR_I[20]), .C(n41266), 
         .D(SHAREDBUS_ADR_I[30]), .Z(n32322)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_871.init = 16'hfffe;
    LUT4 i1_2_lut_adj_872 (.A(\SHAREDBUS_ADR_I[23] ), .B(SHAREDBUS_ADR_I[16]), 
         .Z(n32304)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_adj_872.init = 16'heeee;
    LUT4 i1_4_lut_adj_873 (.A(n32788), .B(n41210), .C(n15), .D(n35884), 
         .Z(FIFOwb_en)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_873.init = 16'h0008;
    LUT4 i1_4_lut_adj_874 (.A(n32774), .B(n41225), .C(n19), .D(n41235), 
         .Z(n32788)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_874.init = 16'h0002;
    LUT4 i30722_4_lut (.A(n35761), .B(n33846), .C(n35739), .D(n41259), 
         .Z(n35884)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30722_4_lut.init = 16'hfffe;
    LUT4 i11_3_lut_adj_875 (.A(ebrEBR_DAT_O[12]), .B(\genblk1.write_data_d [12]), 
         .C(\genblk1.raw_hazard ), .Z(n9_adj_6355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i11_3_lut_adj_875.init = 16'hcaca;
    LUT4 mux_66_i1_4_lut (.A(read_ack), .B(GPIOGPIO_ACK_O), .C(n41180), 
         .D(write_ack), .Z(n1030[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(553[1] 556[2])
    defparam mux_66_i1_4_lut.init = 16'hcfca;
    LUT4 i33240_4_lut (.A(n41194), .B(n41181), .C(n41195), .D(n36343), 
         .Z(n36351)) /* synthesis lut_function=(((C (D))+!B)+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(549[1] 556[2])
    defparam i33240_4_lut.init = 16'hf777;
    LUT4 i1_4_lut_adj_876 (.A(n34104), .B(n41210), .C(n34372), .D(n34444), 
         .Z(n34112)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_876.init = 16'hfffb;
    LUT4 i1_4_lut_adj_877 (.A(n15), .B(n34078), .C(n34396), .D(n34236), 
         .Z(n34104)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_877.init = 16'hfffe;
    LUT4 i1_2_lut_rep_849 (.A(SHAREDBUS_ADR_I[27]), .B(\SHAREDBUS_ADR_I[23] ), 
         .Z(n41254)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_rep_849.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_878 (.A(SHAREDBUS_ADR_I[27]), .B(\SHAREDBUS_ADR_I[23] ), 
         .C(SHAREDBUS_ADR_I[25]), .D(SHAREDBUS_ADR_I[26]), .Z(n32690)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_3_lut_4_lut_adj_878.init = 16'hfffe;
    LUT4 i1_2_lut_adj_879 (.A(SHAREDBUS_ADR_I[20]), .B(reg_04[0]), .Z(n34078)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_adj_879.init = 16'heeee;
    LUT4 i1_2_lut_adj_880 (.A(SHAREDBUS_ADR_I[26]), .B(SHAREDBUS_ADR_I[18]), 
         .Z(n34236)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_adj_880.init = 16'heeee;
    LUT4 i1_4_lut_adj_881 (.A(n41267), .B(n19), .C(n34242), .D(n41276), 
         .Z(n34444)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_881.init = 16'hfffe;
    LUT4 i1_4_lut_adj_882 (.A(n33990), .B(n41210), .C(n34372), .D(n34444), 
         .Z(n33998)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_882.init = 16'hfffb;
    LUT4 i1_4_lut_adj_883 (.A(n15), .B(n33964), .C(n34396), .D(n34236), 
         .Z(n33990)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_883.init = 16'hfffe;
    LUT4 i1_2_lut_adj_884 (.A(SHAREDBUS_ADR_I[20]), .B(reg_04[2]), .Z(n33964)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_adj_884.init = 16'heeee;
    LUT4 i1_4_lut_adj_885 (.A(n34066), .B(n41210), .C(n34372), .D(n34444), 
         .Z(n34074)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_885.init = 16'hfffb;
    LUT4 i1_4_lut_adj_886 (.A(n15), .B(n34040), .C(n34396), .D(n34236), 
         .Z(n34066)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_886.init = 16'hfffe;
    LUT4 i1_2_lut_adj_887 (.A(SHAREDBUS_ADR_I[20]), .B(reg_04[3]), .Z(n34040)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_adj_887.init = 16'heeee;
    LUT4 i1_4_lut_adj_888 (.A(n35910), .B(n41210), .C(n35633), .D(n32980), 
         .Z(n32990)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_888.init = 16'h0400;
    LUT4 i30748_4_lut (.A(n41235), .B(n19), .C(n35808), .D(n35649), 
         .Z(n35910)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30748_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_889 (.A(n34446), .B(n41210), .C(n34372), .D(n34444), 
         .Z(n34454)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_889.init = 16'hfffb;
    LUT4 i1_4_lut_adj_890 (.A(n15), .B(n34420), .C(n34396), .D(n34236), 
         .Z(n34446)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_890.init = 16'hfffe;
    LUT4 i1_2_lut_adj_891 (.A(SHAREDBUS_ADR_I[20]), .B(reg_04[6]), .Z(n34420)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_adj_891.init = 16'heeee;
    LUT4 i1_4_lut_adj_892 (.A(n34142), .B(n41210), .C(n34372), .D(n34444), 
         .Z(n34150)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_892.init = 16'hfffb;
    LUT4 i1_4_lut_adj_893 (.A(n15), .B(n34116), .C(n34396), .D(n34236), 
         .Z(n34142)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_893.init = 16'hfffe;
    LUT4 i1_2_lut_adj_894 (.A(SHAREDBUS_ADR_I[20]), .B(reg_04[7]), .Z(n34116)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_adj_894.init = 16'heeee;
    LUT4 i1_4_lut_adj_895 (.A(n35910), .B(n41210), .C(n35633), .D(n32940), 
         .Z(n32950)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_895.init = 16'h0400;
    LUT4 i1_4_lut_adj_896 (.A(n32028), .B(n19), .C(n41301), .D(SHAREDBUS_ADR_I[24]), 
         .Z(n32038)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_896.init = 16'hfffe;
    LUT4 i1_4_lut_adj_897 (.A(n35761), .B(n32032), .C(\SHAREDBUS_ADR_I[22] ), 
         .D(\SHAREDBUS_ADR_I[23] ), .Z(n32036)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_897.init = 16'hfffe;
    LUT4 i1_2_lut_rep_854 (.A(\SHAREDBUS_ADR_I[23] ), .B(SHAREDBUS_ADR_I[24]), 
         .Z(n41259)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_rep_854.init = 16'heeee;
    LUT4 i30565_2_lut_3_lut_4_lut (.A(\SHAREDBUS_ADR_I[23] ), .B(SHAREDBUS_ADR_I[24]), 
         .C(SHAREDBUS_ADR_I[25]), .D(SHAREDBUS_ADR_I[30]), .Z(n35724)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i30565_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut_adj_898 (.A(n41310), .B(n41301), .C(n41303), .D(n41304), 
         .Z(n35184)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_898.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_899 (.A(n41310), .B(n41301), .C(n41344), 
         .D(n41345), .Z(n34816)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_899.init = 16'h8000;
    LUT4 i1_3_lut_4_lut_adj_900 (.A(n41310), .B(n41301), .C(n41303), .D(SHAREDBUS_ADR_I[30]), 
         .Z(n32774)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_900.init = 16'h0008;
    LUT4 i1_3_lut_4_lut_adj_901 (.A(n41303), .B(\SHAREDBUS_ADR_I[23] ), 
         .C(n33846), .D(n41276), .Z(n33864)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_3_lut_4_lut_adj_901.init = 16'hfffe;
    LUT4 i1_2_lut_rep_859 (.A(SHAREDBUS_ADR_I[30]), .B(\SHAREDBUS_ADR_I[22] ), 
         .Z(n41264)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_rep_859.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut_adj_902 (.A(SHAREDBUS_ADR_I[30]), .B(\SHAREDBUS_ADR_I[22] ), 
         .C(SHAREDBUS_ADR_I[24]), .D(\SHAREDBUS_ADR_I[23] ), .Z(n34396)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_3_lut_4_lut_adj_902.init = 16'hfffe;
    LUT4 i1_2_lut_rep_860 (.A(SHAREDBUS_ADR_I[18]), .B(SHAREDBUS_ADR_I[24]), 
         .Z(n41265)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_rep_860.init = 16'heeee;
    LUT4 i1_2_lut_rep_861 (.A(\SHAREDBUS_ADR_I[29] ), .B(SHAREDBUS_ADR_I[26]), 
         .Z(n41266)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_rep_861.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_903 (.A(\SHAREDBUS_ADR_I[29] ), .B(SHAREDBUS_ADR_I[26]), 
         .C(SHAREDBUS_ADR_I[20]), .D(SHAREDBUS_ADR_I[25]), .Z(n32890)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_3_lut_4_lut_adj_903.init = 16'hfffe;
    LUT4 i1_2_lut_rep_862 (.A(SHAREDBUS_ADR_I[27]), .B(SHAREDBUS_ADR_I[25]), 
         .Z(n41267)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_rep_862.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut_adj_904 (.A(SHAREDBUS_ADR_I[27]), .B(SHAREDBUS_ADR_I[25]), 
         .C(SHAREDBUS_ADR_I[24]), .D(SHAREDBUS_ADR_I[18]), .Z(n32318)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_3_lut_4_lut_adj_904.init = 16'hfffe;
    LUT4 i1_2_lut_rep_863 (.A(\SHAREDBUS_ADR_I[22] ), .B(SHAREDBUS_ADR_I[16]), 
         .Z(n41268)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_rep_863.init = 16'heeee;
    LUT4 i1_2_lut_rep_864 (.A(\SHAREDBUS_ADR_I[23] ), .B(SHAREDBUS_ADR_I[30]), 
         .Z(n41269)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_rep_864.init = 16'heeee;
    LUT4 i30433_2_lut_3_lut_4_lut (.A(\SHAREDBUS_ADR_I[23] ), .B(SHAREDBUS_ADR_I[30]), 
         .C(SHAREDBUS_ADR_I[25]), .D(SHAREDBUS_ADR_I[24]), .Z(n35577)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i30433_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i30692_3_lut_4_lut (.A(\SHAREDBUS_ADR_I[23] ), .B(SHAREDBUS_ADR_I[30]), 
         .C(SHAREDBUS_ADR_I[26]), .D(n19), .Z(n35854)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i30692_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_865 (.A(SHAREDBUS_ADR_I[20]), .B(SHAREDBUS_ADR_I[18]), 
         .Z(n41270)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_rep_865.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_905 (.A(SHAREDBUS_ADR_I[20]), .B(SHAREDBUS_ADR_I[18]), 
         .C(SHAREDBUS_ADR_I[24]), .D(SHAREDBUS_ADR_I[26]), .Z(n32192)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_3_lut_4_lut_adj_905.init = 16'hfffe;
    LUT4 i1_2_lut_rep_871 (.A(SHAREDBUS_ADR_I[16]), .B(\SHAREDBUS_ADR_I[29] ), 
         .Z(n41276)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_rep_871.init = 16'heeee;
    LUT4 i1_2_lut_rep_815_3_lut_4_lut (.A(SHAREDBUS_ADR_I[16]), .B(\SHAREDBUS_ADR_I[29] ), 
         .C(\SHAREDBUS_ADR_I[22] ), .D(SHAREDBUS_ADR_I[20]), .Z(n41220)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_rep_815_3_lut_4_lut.init = 16'hfffe;
    LUT4 i30553_2_lut_3_lut_4_lut (.A(SHAREDBUS_ADR_I[16]), .B(\SHAREDBUS_ADR_I[29] ), 
         .C(SHAREDBUS_ADR_I[26]), .D(SHAREDBUS_ADR_I[20]), .Z(n35712)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i30553_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i30601_2_lut (.A(SHAREDBUS_ADR_I[26]), .B(SHAREDBUS_ADR_I[27]), 
         .Z(n35761)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i30601_2_lut.init = 16'heeee;
    LUT4 i12_3_lut_adj_906 (.A(n9_adj_6452), .B(\genblk1.EBR_DAT_I_d [16]), 
         .C(\genblk1.EBR_SEL_I_d [2]), .Z(\genblk1.write_data_23__N_3549 [0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i12_3_lut_adj_906.init = 16'hcaca;
    LUT4 i1_4_lut_adj_907 (.A(n35910), .B(n41210), .C(n35633), .D(n33100), 
         .Z(n33110)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_907.init = 16'h0400;
    LUT4 i1_3_lut_adj_908 (.A(n41300), .B(n29), .C(n41299), .Z(n15)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_3_lut_adj_908.init = 16'hfefe;
    LUT4 i1_4_lut_4_lut (.A(n41310), .B(n33954), .C(REF_CLK_c_enable_424), 
         .D(n30231), .Z(n31183)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_4_lut_4_lut.init = 16'h4000;
    LUT4 i1_4_lut_4_lut_adj_909 (.A(n41310), .B(n33332), .C(n41246), .D(n35577), 
         .Z(n33356)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_4_lut_4_lut_adj_909.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_adj_910 (.A(n41310), .B(n19), .C(n32814), .D(n41210), 
         .Z(n32828)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(797[20:79])
    defparam i1_4_lut_4_lut_adj_910.init = 16'hfdff;
    PFUMX i23 (.BLUT(n8_c), .ALUT(n11_adj_6446), .C0(n37907), .Z(SHAREDBUS_DAT_O[8]));
    PFUMX i23_adj_911 (.BLUT(n8_adj_6454), .ALUT(n11_adj_6444), .C0(n37909), 
          .Z(SHAREDBUS_DAT_O[27]));
    PFUMX i23_adj_912 (.BLUT(n8_adj_6455), .ALUT(n11_adj_6442), .C0(n37910), 
          .Z(SHAREDBUS_DAT_O[20]));
    PFUMX i23_adj_913 (.BLUT(n8_adj_6456), .ALUT(n11_adj_6440), .C0(n37911), 
          .Z(SHAREDBUS_DAT_O[19]));
    PFUMX i23_adj_914 (.BLUT(n8_adj_6457), .ALUT(n11_adj_6438), .C0(n37909), 
          .Z(SHAREDBUS_DAT_O[26]));
    PFUMX i23_adj_915 (.BLUT(n8_adj_6458), .ALUT(n11_adj_6436), .C0(n37911), 
          .Z(SHAREDBUS_DAT_O[16]));
    PFUMX i23_adj_916 (.BLUT(n8_adj_6459), .ALUT(n11_adj_6434), .C0(n37908), 
          .Z(SHAREDBUS_DAT_O[31]));
    PFUMX i23_adj_917 (.BLUT(n8_adj_6460), .ALUT(n11_adj_6432), .C0(n37908), 
          .Z(SHAREDBUS_DAT_O[30]));
    PFUMX i23_adj_918 (.BLUT(n8_adj_6461), .ALUT(n11_adj_6430), .C0(n37907), 
          .Z(SHAREDBUS_DAT_O[5]));
    PFUMX i23_adj_919 (.BLUT(n8_adj_6462), .ALUT(n11_adj_6429), .C0(n37912), 
          .Z(SHAREDBUS_DAT_O[12]));
    PFUMX i23_adj_920 (.BLUT(n8_adj_6463), .ALUT(n11_adj_6427), .C0(n37910), 
          .Z(SHAREDBUS_DAT_O[23]));
    PFUMX i23_adj_921 (.BLUT(n8_adj_6464), .ALUT(n11_adj_6426), .C0(n37907), 
          .Z(SHAREDBUS_DAT_O[1]));
    PFUMX i23_adj_922 (.BLUT(n8_adj_6465), .ALUT(n11_adj_6425), .C0(n37913), 
          .Z(SHAREDBUS_DAT_O[10]));
    PFUMX i23_adj_923 (.BLUT(n8_adj_6466), .ALUT(n11_adj_6423), .C0(n37907), 
          .Z(SHAREDBUS_DAT_O[0]));
    PFUMX i23_adj_924 (.BLUT(n8_adj_6467), .ALUT(n11_adj_6422), .C0(n37913), 
          .Z(SHAREDBUS_DAT_O[7]));
    PFUMX i23_adj_925 (.BLUT(n8_adj_6468), .ALUT(n11_adj_6420), .C0(n37910), 
          .Z(SHAREDBUS_DAT_O[22]));
    PFUMX i23_adj_926 (.BLUT(n8_adj_6469), .ALUT(n11_adj_6418), .C0(n41194), 
          .Z(SHAREDBUS_DAT_O[6]));
    PFUMX i23_adj_927 (.BLUT(n8_adj_6470), .ALUT(n11_adj_6416), .C0(n41194), 
          .Z(SHAREDBUS_DAT_O[4]));
    PFUMX i21 (.BLUT(n3_adj_6471), .ALUT(n9_adj_6414), .C0(n37908), .Z(SHAREDBUS_DAT_O[28]));
    PFUMX i23_adj_928 (.BLUT(n8_adj_6472), .ALUT(n11_adj_6412), .C0(n41194), 
          .Z(SHAREDBUS_DAT_O[3]));
    PFUMX i23_adj_929 (.BLUT(n8_adj_6473), .ALUT(n11_adj_6410), .C0(n41194), 
          .Z(SHAREDBUS_DAT_O[2]));
    PFUMX i21_adj_930 (.BLUT(n3_adj_6474), .ALUT(n9_adj_6408), .C0(n37910), 
          .Z(SHAREDBUS_DAT_O[21]));
    LUT4 i1_4_lut_adj_931 (.A(n35910), .B(n41210), .C(n35633), .D(n33060), 
         .Z(n33070)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_931.init = 16'h0400;
    PFUMX i21_adj_932 (.BLUT(n3_adj_6475), .ALUT(n9_adj_6406), .C0(n37909), 
          .Z(SHAREDBUS_DAT_O[25]));
    PFUMX i21_adj_933 (.BLUT(n3_adj_6476), .ALUT(n9_adj_6404), .C0(n37911), 
          .Z(SHAREDBUS_DAT_O[18]));
    PFUMX i23_adj_934 (.BLUT(n8_adj_6477), .ALUT(n11_adj_6402), .C0(n37911), 
          .Z(SHAREDBUS_DAT_O[17]));
    LUT4 i15_4_lut (.A(n33368), .B(reg_00[24]), .C(n41185), .D(n33214), 
         .Z(n21)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(89[9:19])
    defparam i15_4_lut.init = 16'hcac0;
    PFUMX i30 (.BLUT(n3_adj_6478), .ALUT(n14_adj_6398), .C0(n37912), .Z(SHAREDBUS_DAT_O[15]));
    PFUMX i23_adj_935 (.BLUT(n8_adj_6479), .ALUT(n11_adj_6396), .C0(n37912), 
          .Z(SHAREDBUS_DAT_O[14]));
    PFUMX i30_adj_936 (.BLUT(n3_adj_6480), .ALUT(n14_adj_6394), .C0(n37912), 
          .Z(SHAREDBUS_DAT_O[13]));
    PFUMX i23_adj_937 (.BLUT(n8_adj_6481), .ALUT(n11_adj_6392), .C0(n37908), 
          .Z(SHAREDBUS_DAT_O[29]));
    PFUMX i30_adj_938 (.BLUT(n3_adj_6482), .ALUT(n14_adj_6391), .C0(n37913), 
          .Z(SHAREDBUS_DAT_O[11]));
    PFUMX i30_adj_939 (.BLUT(n3_adj_6483), .ALUT(n14), .C0(n37913), .Z(SHAREDBUS_DAT_O[9]));
    PFUMX i30_adj_940 (.BLUT(n11_adj_6484), .ALUT(n14_adj_6485), .C0(n37909), 
          .Z(SHAREDBUS_DAT_O[24]));
    LUT4 i1_4_lut_adj_941 (.A(n35910), .B(n41210), .C(n35633), .D(n32864), 
         .Z(n32874)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_941.init = 16'h0400;
    PFUMX i9 (.BLUT(n13_adj_6486), .ALUT(n17_adj_6388), .C0(n37931), .Z(n19_adj_6487));
    PFUMX i9_adj_942 (.BLUT(n13_adj_6488), .ALUT(n17_adj_6387), .C0(n37931), 
          .Z(n19_adj_6489));
    PFUMX i9_adj_943 (.BLUT(n13_adj_6490), .ALUT(n17_adj_6386), .C0(n37931), 
          .Z(n19_adj_6491));
    PFUMX i9_adj_944 (.BLUT(n13_adj_6492), .ALUT(n17_adj_6385), .C0(n37930), 
          .Z(n19_adj_6493));
    LUT4 i1_4_lut_adj_945 (.A(\SHAREDBUS_ADR_I[5] ), .B(n41346), .C(n33948), 
         .D(\SHAREDBUS_ADR_I[7] ), .Z(n33954)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_945.init = 16'h1000;
    PFUMX i9_adj_946 (.BLUT(n11_adj_6494), .ALUT(n15_adj_6384), .C0(n37929), 
          .Z(n17_adj_6495));
    PFUMX i9_adj_947 (.BLUT(n13_adj_6496), .ALUT(n17_adj_6383), .C0(n37929), 
          .Z(n19_adj_6497));
    PFUMX i9_adj_948 (.BLUT(n13_adj_6498), .ALUT(n17_adj_6382), .C0(n37928), 
          .Z(n19_adj_6499));
    PFUMX i9_adj_949 (.BLUT(n13_adj_6500), .ALUT(n17_adj_6381), .C0(n37928), 
          .Z(n19_adj_6501));
    PFUMX i9_adj_950 (.BLUT(n13_adj_6502), .ALUT(n17_adj_6380), .C0(n37927), 
          .Z(n19_adj_6503));
    PFUMX i14 (.BLUT(n9_adj_6504), .ALUT(n17_adj_6379), .C0(n37927), .Z(n19_adj_6505));
    PFUMX mux_108_i9 (.BLUT(GPOwb_DAT_O[8]), .ALUT(n295[8]), .C0(n37926), 
          .Z(n328[8])) /* synthesis LSE_LINE_FILE_ID=60, LSE_LCOL=13, LSE_RCOL=22, LSE_LLINE=54, LSE_RLINE=54 */ ;
    PFUMX mux_108_i6 (.BLUT(GPOwb_DAT_O[5]), .ALUT(n295[5]), .C0(n37926), 
          .Z(n328[5])) /* synthesis LSE_LINE_FILE_ID=60, LSE_LCOL=13, LSE_RCOL=22, LSE_LLINE=54, LSE_RLINE=54 */ ;
    PFUMX mux_108_i2 (.BLUT(GPOwb_DAT_O[1]), .ALUT(n295[1]), .C0(n37926), 
          .Z(n328[1])) /* synthesis LSE_LINE_FILE_ID=60, LSE_LCOL=13, LSE_RCOL=22, LSE_LLINE=54, LSE_RLINE=54 */ ;
    PFUMX mux_8_i1 (.BLUT(n1063[0]), .ALUT(SHAREDBUS_ACK_O_N_91[0]), .C0(n36351), 
          .Z(n949[0])) /* synthesis LSE_LINE_FILE_ID=60, LSE_LCOL=13, LSE_RCOL=22, LSE_LLINE=54, LSE_RLINE=54 */ ;
    LUT4 i1_2_lut_adj_951 (.A(n954[0]), .B(PIO_DATAI[0]), .Z(n33948)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_951.init = 16'h8888;
    PFUMX mux_108_i1 (.BLUT(GPOwb_DAT_O[0]), .ALUT(n295[0]), .C0(n37926), 
          .Z(n328[0])) /* synthesis LSE_LINE_FILE_ID=60, LSE_LCOL=13, LSE_RCOL=22, LSE_LLINE=54, LSE_RLINE=54 */ ;
    PFUMX i13827 (.BLUT(n4_adj_6377), .ALUT(n6_adj_6376), .C0(n41189), 
          .Z(n8_adj_6506));
    PFUMX i13795 (.BLUT(n4_adj_6375), .ALUT(n6_adj_6374), .C0(n37932), 
          .Z(n8_adj_6507));
    PFUMX i9_adj_952 (.BLUT(n11_adj_6373), .ALUT(n15_adj_6372), .C0(n37932), 
          .Z(n17_adj_6508));
    PFUMX i13687 (.BLUT(n4_adj_6371), .ALUT(n6_adj_6370), .C0(n37932), 
          .Z(n8_adj_6509));
    PFUMX i13655 (.BLUT(n4), .ALUT(n6), .C0(n37932), .Z(n8_adj_6510));
    PFUMX i9_adj_953 (.BLUT(n13_adj_6369), .ALUT(n17_adj_6368), .C0(n37931), 
          .Z(n19_adj_6511));
    PFUMX i9_adj_954 (.BLUT(n13_adj_6367), .ALUT(n17_adj_6366), .C0(n37930), 
          .Z(n19_adj_6512));
    PFUMX i9_adj_955 (.BLUT(n13_adj_6365), .ALUT(n17_adj_6364), .C0(n37929), 
          .Z(n19_adj_6513));
    PFUMX i14_adj_956 (.BLUT(n15_adj_6363), .ALUT(n3_adj_6362), .C0(n37930), 
          .Z(n16_adj_6514));
    PFUMX i14_adj_957 (.BLUT(n15_adj_6361), .ALUT(n3_adj_6360), .C0(n37929), 
          .Z(n16_adj_6515));
    PFUMX i9_adj_958 (.BLUT(n13), .ALUT(n17), .C0(n37927), .Z(n19_adj_6516));
    PFUMX i14_adj_959 (.BLUT(n15_adj_6359), .ALUT(n3_adj_6358), .C0(n37930), 
          .Z(n16_adj_6517));
    PFUMX i14_adj_960 (.BLUT(n15_adj_6357), .ALUT(n3_adj_6356), .C0(n37928), 
          .Z(n16_adj_6518));
    LUT4 i1_4_lut_adj_961 (.A(n34180), .B(n41210), .C(n34372), .D(n34444), 
         .Z(n34188)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_961.init = 16'hfffb;
    LUT4 i1_4_lut_adj_962 (.A(n15), .B(n34154), .C(n34396), .D(n34236), 
         .Z(n34180)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_962.init = 16'hfffe;
    PFUMX i31 (.BLUT(n15_adj_6354), .ALUT(n3_adj_6353), .C0(n41189), .Z(n16_adj_6519));
    PFUMX i31_adj_963 (.BLUT(n15_adj_6352), .ALUT(n3_adj_6351), .C0(n41189), 
          .Z(n16_adj_6520));
    LUT4 i1_2_lut_adj_964 (.A(SHAREDBUS_ADR_I[20]), .B(reg_04[18]), .Z(n34154)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_adj_964.init = 16'heeee;
    PFUMX i31_adj_965 (.BLUT(n15_adj_6350), .ALUT(n3_adj_6349), .C0(n37927), 
          .Z(n16_adj_6521));
    PFUMX i31_adj_966 (.BLUT(n15_adj_6348), .ALUT(n3_adj_6347), .C0(n37928), 
          .Z(n16_adj_6522));
    LUT4 i1_4_lut_adj_967 (.A(n34028), .B(n41210), .C(n34372), .D(n34444), 
         .Z(n34036)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_967.init = 16'hfffb;
    LUT4 i1_4_lut_adj_968 (.A(n15), .B(n34002), .C(n34396), .D(n34236), 
         .Z(n34028)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_968.init = 16'hfffe;
    LUT4 i1_2_lut_adj_969 (.A(SHAREDBUS_ADR_I[20]), .B(reg_04[25]), .Z(n34002)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_adj_969.init = 16'heeee;
    LUT4 i1_4_lut_adj_970 (.A(n35910), .B(n41210), .C(n35633), .D(n33020), 
         .Z(n33030)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_970.init = 16'h0400;
    LUT4 i1_4_lut_adj_971 (.A(n34256), .B(n41210), .C(n34372), .D(n34444), 
         .Z(n34264)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_971.init = 16'hfffb;
    LUT4 i1_4_lut_adj_972 (.A(n15), .B(n34230), .C(n34396), .D(n34236), 
         .Z(n34256)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_972.init = 16'hfffe;
    LUT4 i1_2_lut_adj_973 (.A(SHAREDBUS_ADR_I[20]), .B(reg_04[21]), .Z(n34230)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_adj_973.init = 16'heeee;
    LUT4 i1_4_lut_adj_974 (.A(n34332), .B(n41210), .C(n34372), .D(n34444), 
         .Z(n34340)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_974.init = 16'hfffb;
    LUT4 i1_4_lut_adj_975 (.A(n15), .B(n34306), .C(n34396), .D(n34236), 
         .Z(n34332)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_975.init = 16'hfffe;
    LUT4 i1_2_lut_adj_976 (.A(SHAREDBUS_ADR_I[20]), .B(reg_04[28]), .Z(n34306)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_adj_976.init = 16'heeee;
    LUT4 i1_4_lut_adj_977 (.A(n34408), .B(n41210), .C(n34372), .D(n34444), 
         .Z(n34416)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_977.init = 16'hfffb;
    LUT4 i1_4_lut_adj_978 (.A(n15), .B(n34382), .C(n34396), .D(n34236), 
         .Z(n34408)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_978.init = 16'hfffe;
    LUT4 i1_2_lut_adj_979 (.A(SHAREDBUS_ADR_I[20]), .B(reg_04[15]), .Z(n34382)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_adj_979.init = 16'heeee;
    LUT4 i1_4_lut_adj_980 (.A(n34370), .B(n41210), .C(n34372), .D(n34444), 
         .Z(n34378)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_980.init = 16'hfffb;
    LUT4 i1_4_lut_adj_981 (.A(n15), .B(n34344), .C(n34396), .D(n34236), 
         .Z(n34370)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_981.init = 16'hfffe;
    LUT4 i1_2_lut_adj_982 (.A(SHAREDBUS_ADR_I[20]), .B(reg_04[13]), .Z(n34344)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_adj_982.init = 16'heeee;
    LUT4 i1_4_lut_adj_983 (.A(n34294), .B(n41210), .C(n34372), .D(n34444), 
         .Z(n34302)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_983.init = 16'hfffb;
    LUT4 i1_4_lut_adj_984 (.A(n15), .B(n34268), .C(n34396), .D(n34236), 
         .Z(n34294)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_984.init = 16'hfffe;
    LUT4 i1_2_lut_adj_985 (.A(SHAREDBUS_ADR_I[20]), .B(reg_04[11]), .Z(n34268)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_adj_985.init = 16'heeee;
    LUT4 i10_3_lut_adj_986 (.A(ebrEBR_DAT_O[11]), .B(\genblk1.write_data_d [11]), 
         .C(\genblk1.raw_hazard ), .Z(n11_adj_6346)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(247[11:21])
    defparam i10_3_lut_adj_986.init = 16'hcaca;
    LUT4 i1_4_lut_adj_987 (.A(n34218), .B(n41210), .C(n34372), .D(n34444), 
         .Z(n34226)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_987.init = 16'hfffb;
    LUT4 i1_4_lut_adj_988 (.A(n15), .B(n34192), .C(n34396), .D(n34236), 
         .Z(n34218)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_4_lut_adj_988.init = 16'hfffe;
    LUT4 i1_2_lut_adj_989 (.A(SHAREDBUS_ADR_I[20]), .B(reg_04[9]), .Z(n34192)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(661[20:70])
    defparam i1_2_lut_adj_989.init = 16'heeee;
    LUT4 i1_4_lut_adj_990 (.A(n32074), .B(n35930), .C(n41225), .D(n19), 
         .Z(n32084)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_990.init = 16'h0002;
    LUT4 i1_4_lut_adj_991 (.A(SHAREDBUS_ADR_I[30]), .B(n41268), .C(n41303), 
         .D(n32054), .Z(n32074)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_991.init = 16'h0100;
    LUT4 i30768_4_lut (.A(n15), .B(n35761), .C(n35866), .D(n41242), 
         .Z(n35930)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30768_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_992 (.A(n41301), .B(n41310), .C(write_ack_adj_6523), 
         .D(read_ack_adj_6524), .Z(n32054)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_992.init = 16'h8880;
    \spi(SLAVE_NUMBER=32'b01,CLKCNT_WIDTH=16)  spi (.sclk_N_5010(sclk_N_5010), 
            .IO_SCK_c(IO_SCK_c), .spiSPI_ACK_O(spiSPI_ACK_O), .REF_CLK_c(REF_CLK_c), 
            .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), .spiSPI_DAT_O({spiSPI_DAT_O}), 
            .rx_shift_data_31__N_4339(rx_shift_data_31__N_4339), .n41328(n41328), 
            .dw10_cs_N_4471(dw10_cs_N_4471), .REF_CLK_c_enable_1453(REF_CLK_c_enable_1453), 
            .IO_MISO_c(IO_MISO_c), .dw00_cs_N_4467(dw00_cs_N_4467), .IO_0_c_0(IO_0_c_0), 
            .GND_net(GND_net), .VCC_net(VCC_net), .IO_MOSI_c(IO_MOSI_c), 
            .n41329(n41329), .n41330(n41330), .n41331(n41331), .n41332(n41332), 
            .n41333(n41333), .n41334(n41334), .n41335(n41335), .\SHAREDBUS_DAT_I[8] (\SHAREDBUS_DAT_I[8] ), 
            .\SHAREDBUS_DAT_I[9] (\SHAREDBUS_DAT_I[9] ), .\SHAREDBUS_DAT_I[10] (\SHAREDBUS_DAT_I[10] ), 
            .\SHAREDBUS_DAT_I[11] (\SHAREDBUS_DAT_I[11] ), .\SHAREDBUS_DAT_I[12] (\SHAREDBUS_DAT_I[12] ), 
            .\SHAREDBUS_DAT_I[13] (\SHAREDBUS_DAT_I[13] ), .\SHAREDBUS_DAT_I[14] (\SHAREDBUS_DAT_I[14] ), 
            .\SHAREDBUS_DAT_I[15] (\SHAREDBUS_DAT_I[15] ), .n41336(n41336), 
            .n41337(n41337), .n41338(n41338), .n41339(n41339), .n41340(n41340), 
            .n41341(n41341), .n41342(n41342), .n41343(n41343), .\SHAREDBUS_DAT_I[24] (\SHAREDBUS_DAT_I[24] ), 
            .\SHAREDBUS_DAT_I[25] (\SHAREDBUS_DAT_I[25] ), .\SHAREDBUS_DAT_I[26] (\SHAREDBUS_DAT_I[26] ), 
            .\SHAREDBUS_DAT_I[27] (\SHAREDBUS_DAT_I[27] ), .\SHAREDBUS_DAT_I[28] (\SHAREDBUS_DAT_I[28] ), 
            .\SHAREDBUS_DAT_I[29] (\SHAREDBUS_DAT_I[29] ), .\SHAREDBUS_DAT_I[30] (\SHAREDBUS_DAT_I[30] ), 
            .\SHAREDBUS_DAT_I[31] (\SHAREDBUS_DAT_I[31] ), .n45179(n45179), 
            .n41225(n41225), .\LM32D_ADR_O[1] (LM32D_ADR_O[1]), .n41380(n41380), 
            .\LM32D_ADR_O[0] (LM32D_ADR_O[0]), .n30156(n30156), .n41246(n41246), 
            .n30986(n30986), .n41310(n41310), .n41304(n41304), .n35042(n35042), 
            .\inst_reg[15] (\inst_reg[15] ), .n10865(n10865), .n41191(n41191), 
            .n41345(n41345), .n41344(n41344), .n41347(n41347), .n34742(n34742), 
            .SPI_INT_O_N_4422(SPI_INT_O_N_4422), .SPI_INT_O_N_4417(SPI_INT_O_N_4417), 
            .SPI_INT_O_N_4421(SPI_INT_O_N_4421), .n953({n953}), .n954({n954}), 
            .n34304(n34304), .\genblk1.wait_one_tick_done (\genblk1.wait_one_tick_done )) /* synthesis syn_module_defined=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(771[2] 790[34])
    \wb_ebr_ctrl(SIZE=32768)  ebr (.\genblk1.write_data_7__N_3573 ({\genblk1.write_data_7__N_3573 }), 
            .REF_CLK_c(REF_CLK_c), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .n41324(n41324), .VCC_net(VCC_net), .ebrEBR_DAT_O({ebrEBR_DAT_O}), 
            .\genblk1.read_address[10] (\genblk1.read_address[10] ), .\genblk1.write_address[10] (\genblk1.write_address[10] ), 
            .n3700(n3700), .n5386(n5386), .n5085(n5085), .n41345(n41345), 
            .n3432(n3432), .n41323(n41323), .n41255(n41255), .\genblk1.state[2] (\genblk1.state[2] ), 
            .GND_net(GND_net), .\genblk1.raw_hazard (\genblk1.raw_hazard ), 
            .ebrEBR_ACK_O(ebrEBR_ACK_O), .\genblk1.write_data_23__N_3541 ({\genblk1.write_data_23__N_3541 }), 
            .\genblk1.write_data_23__N_3549 ({Open_1, Open_2, Open_3, 
            Open_4, Open_5, Open_6, Open_7, \genblk1.write_data_23__N_3549 [0]}), 
            .\genblk1.write_data_31__N_3525 ({\genblk1.write_data_31__N_3525 }), 
            .\genblk1.write_data_15__N_3557 ({\genblk1.write_data_15__N_3557 }), 
            .n12390(n12390), .LM32D_DAT_O({LM32D_DAT_O}), .\genblk1.read_data[20] (\genblk1.read_data [20]), 
            .\genblk1.EBR_SEL_I_d[2] (\genblk1.EBR_SEL_I_d [2]), .\genblk1.EBR_DAT_I_d[9] (\genblk1.EBR_DAT_I_d [9]), 
            .\genblk1.EBR_DAT_I_d[10] (\genblk1.EBR_DAT_I_d [10]), .\genblk1.EBR_DAT_I_d[11] (\genblk1.EBR_DAT_I_d [11]), 
            .\genblk1.EBR_DAT_I_d[12] (\genblk1.EBR_DAT_I_d [12]), .\genblk1.EBR_DAT_I_d[13] (\genblk1.EBR_DAT_I_d [13]), 
            .\genblk1.EBR_DAT_I_d[14] (\genblk1.EBR_DAT_I_d [14]), .\genblk1.EBR_DAT_I_d[15] (\genblk1.EBR_DAT_I_d [15]), 
            .\genblk1.EBR_DAT_I_d[16] (\genblk1.EBR_DAT_I_d [16]), .\genblk1.EBR_DAT_I_d[17] (\genblk1.EBR_DAT_I_d [17]), 
            .\genblk1.EBR_DAT_I_d[18] (\genblk1.EBR_DAT_I_d [18]), .\genblk1.EBR_DAT_I_d[19] (\genblk1.EBR_DAT_I_d [19]), 
            .\genblk1.EBR_DAT_I_d[21] (\genblk1.EBR_DAT_I_d [21]), .\genblk1.EBR_DAT_I_d[22] (\genblk1.EBR_DAT_I_d [22]), 
            .\genblk1.EBR_DAT_I_d[23] (\genblk1.EBR_DAT_I_d [23]), .\genblk1.EBR_DAT_I_d[25] (\genblk1.EBR_DAT_I_d [25]), 
            .\genblk1.EBR_DAT_I_d[26] (\genblk1.EBR_DAT_I_d [26]), .\genblk1.EBR_DAT_I_d[27] (\genblk1.EBR_DAT_I_d [27]), 
            .\genblk1.EBR_DAT_I_d[28] (\genblk1.EBR_DAT_I_d [28]), .\genblk1.EBR_DAT_I_d[29] (\genblk1.EBR_DAT_I_d [29]), 
            .\genblk1.EBR_DAT_I_d[30] (\genblk1.EBR_DAT_I_d [30]), .\genblk1.EBR_DAT_I_d[31] (\genblk1.EBR_DAT_I_d [31]), 
            .\genblk1.EBR_SEL_I_d[1] (\genblk1.EBR_SEL_I_d [1]), .n41238(n41238), 
            .n41309(n41309), .\genblk1.EBR_SEL_I_d[3] (\genblk1.EBR_SEL_I_d [3]), 
            .n41239(n41239), .\genblk1.write_data_d[2] (\genblk1.write_data_d [2]), 
            .\genblk1.write_data_d[3] (\genblk1.write_data_d [3]), .\genblk1.write_data_d[4] (\genblk1.write_data_d [4]), 
            .\genblk1.write_data_d[6] (\genblk1.write_data_d [6]), .\genblk1.write_data_d[7] (\genblk1.write_data_d [7]), 
            .\genblk1.write_data_d[9] (\genblk1.write_data_d [9]), .\genblk1.write_data_d[10] (\genblk1.write_data_d [10]), 
            .\genblk1.write_data_d[11] (\genblk1.write_data_d [11]), .\genblk1.write_data_d[12] (\genblk1.write_data_d [12]), 
            .\genblk1.write_data_d[13] (\genblk1.write_data_d [13]), .\genblk1.write_data_d[14] (\genblk1.write_data_d [14]), 
            .\genblk1.write_data_d[15] (\genblk1.write_data_d [15]), .\genblk1.write_data_d[16] (\genblk1.write_data_d [16]), 
            .\genblk1.write_data_d[17] (\genblk1.write_data_d [17]), .\genblk1.write_data_d[18] (\genblk1.write_data_d [18]), 
            .\genblk1.write_data_d[19] (\genblk1.write_data_d [19]), .\genblk1.write_data_d[20] (\genblk1.write_data_d [20]), 
            .\genblk1.write_data_d[21] (\genblk1.write_data_d [21]), .\genblk1.write_data_d[22] (\genblk1.write_data_d [22]), 
            .\genblk1.write_data_d[23] (\genblk1.write_data_d [23]), .\genblk1.write_data_d[24] (\genblk1.write_data_d [24]), 
            .\genblk1.write_data_d[25] (\genblk1.write_data_d [25]), .\genblk1.write_data_d[26] (\genblk1.write_data_d [26]), 
            .\genblk1.write_data_d[27] (\genblk1.write_data_d [27]), .\genblk1.write_data_d[28] (\genblk1.write_data_d [28]), 
            .\genblk1.write_data_d[29] (\genblk1.write_data_d [29]), .\genblk1.write_data_d[30] (\genblk1.write_data_d [30]), 
            .\genblk1.write_data_d[31] (\genblk1.write_data_d [31]), .n41461(n41461), 
            .n10004(n10004), .\genblk1.pmi_address[3] (\genblk1.pmi_address[3] ), 
            .n10006(n10006), .\genblk1.pmi_address[4] (\genblk1.pmi_address[4] ), 
            .n10008(n10008), .\genblk1.pmi_address[5] (\genblk1.pmi_address[5] ), 
            .n41488(n41488), .\genblk1.pmi_address[6] (\genblk1.pmi_address[6] ), 
            .n10012(n10012), .\genblk1.pmi_address[7] (\genblk1.pmi_address[7] ), 
            .n41485(n41485), .\genblk1.pmi_address[8] (\genblk1.pmi_address[8] ), 
            .n10016(n10016), .\genblk1.pmi_address[9] (\genblk1.pmi_address[9] ), 
            .n10018(n10018), .\genblk1.pmi_address[10] (\genblk1.pmi_address[10] ), 
            .n41482(n41482), .\genblk1.pmi_address[11] (\genblk1.pmi_address[11] ), 
            .n10022(n10022), .\genblk1.pmi_address[12] (\genblk1.pmi_address[12] ), 
            .n10024(n10024), .\genblk1.pmi_address[13] (\genblk1.pmi_address[13] ), 
            .n10026(n10026), .\genblk1.pmi_address[14] (\genblk1.pmi_address[14] ), 
            .n10028(n10028), .n41221(n41221), .n19(n19), .n41304(n41304), 
            .n41321(n41321), .n41195(n41195), .n5(n5_adj_6525), .n35788(n35788), 
            .n41298(n41298), .n20000(n20000), .n41300(n41300), .n41299(n41299), 
            .\SHAREDBUS_ADR_I[10] (\SHAREDBUS_ADR_I[10] ), .n41310(n41310), 
            .n41301(n41301), .\SHAREDBUS_ADR_I[7] (\SHAREDBUS_ADR_I[7] ), 
            .n41346(n41346), .\SHAREDBUS_ADR_I[5] (\SHAREDBUS_ADR_I[5] ), 
            .n41347(n41347), .n41344(n41344), .n6038(n6038), .n15(n15_adj_6526), 
            .n41259(n41259), .n29(n29), .\SHAREDBUS_ADR_I[26] (SHAREDBUS_ADR_I[26]), 
            .\genblk1.read_data[6] (\genblk1.read_data [6]), .n41268(n41268), 
            .n41273(n41273), .n41242(n41242), .n41237(n41237), .\genblk1.read_data[7] (\genblk1.read_data [7]), 
            .n41246(n41246), .\SHAREDBUS_ADR_I[31] (SHAREDBUS_ADR_I[31]), 
            .\SHAREDBUS_ADR_I[15] (SHAREDBUS_ADR_I[15]), .n41222(n41222), 
            .\genblk1.write_data_23__N_3549[7] (\genblk1.write_data_23__N_3549 [7]), 
            .\genblk1.write_data_23__N_3549[6] (\genblk1.write_data_23__N_3549 [6]), 
            .\genblk1.write_data_23__N_3549[5] (\genblk1.write_data_23__N_3549 [5]), 
            .\genblk1.write_data_23__N_3549[3] (\genblk1.write_data_23__N_3549 [3]), 
            .n35840(n35840), .n41260(n41260), .\SHAREDBUS_ADR_I[16] (SHAREDBUS_ADR_I[16]), 
            .\genblk1.write_data_23__N_3549[2] (\genblk1.write_data_23__N_3549 [2]), 
            .n11843(n11843), .\LM32D_ADR_O[1] (LM32D_ADR_O[1]), .n41380(n41380), 
            .n3485(n3485), .n6034(n6034), .n41292(n41292), .n19822(n19822), 
            .n11831(n11831), .n41307(n41307), .n41390(n41390), .n41306(n41306), 
            .n33(n33), .n71(n71), .n3486(n3486), .\counter[2] (\counter[2] ), 
            .n76(n82_adj_325[0]), .n21(n21_adj_6527), .\genblk1.read_data[24] (\genblk1.read_data [24]), 
            .\genblk1.write_data_23__N_3549[1] (\genblk1.write_data_23__N_3549 [1]), 
            .\genblk1.write_data_31__N_3533[7] (\genblk1.write_data_31__N_3533 [7]), 
            .\genblk1.write_data_31__N_3533[6] (\genblk1.write_data_31__N_3533 [6]), 
            .\genblk1.write_data_31__N_3533[5] (\genblk1.write_data_31__N_3533 [5]), 
            .\genblk1.write_data_31__N_3533[4] (\genblk1.write_data_31__N_3533 [4]), 
            .\genblk1.write_data_31__N_3533[3] (\genblk1.write_data_31__N_3533 [3]), 
            .\genblk1.read_data[2] (\genblk1.read_data [2]), .\genblk1.read_data[3] (\genblk1.read_data [3]), 
            .\genblk1.write_data_31__N_3533[2] (\genblk1.write_data_31__N_3533 [2]), 
            .\genblk1.write_data_31__N_3533[1] (\genblk1.write_data_31__N_3533 [1]), 
            .\genblk1.write_data_15__N_3565[7] (\genblk1.write_data_15__N_3565 [7]), 
            .\genblk1.write_data_15__N_3565[6] (\genblk1.write_data_15__N_3565 [6]), 
            .\genblk1.write_data_15__N_3565[5] (\genblk1.write_data_15__N_3565 [5]), 
            .\genblk1.read_data[4] (\genblk1.read_data [4]), .\genblk1.write_data_15__N_3565[4] (\genblk1.write_data_15__N_3565 [4]), 
            .\genblk1.write_data_15__N_3565[3] (\genblk1.write_data_15__N_3565 [3]), 
            .\genblk1.write_data_15__N_3565[2] (\genblk1.write_data_15__N_3565 [2]), 
            .\genblk1.write_data_15__N_3565[1] (\genblk1.write_data_15__N_3565 [1])) /* synthesis syn_module_defined=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(668[2] 682[36])
    arbiter2 arbiter (.LM32D_WE_O(LM32D_WE_O), .n41380(n41380), .n45079(n45079), 
            .n70(n82_adj_325[2]), .n10004(n10004), .n45080(n45080), .n67(n82_adj_325[3]), 
            .n10006(n10006), .n64(n82_adj_325[4]), .n10008(n10008), .n58(n82_adj_325[6]), 
            .n10012(n10012), .n52(n82_adj_325[8]), .n10016(n10016), .n49(n82_adj_325[9]), 
            .n10018(n10018), .n43(n82_adj_325[11]), .n10022(n10022), .n45076(n45076), 
            .n40(n82_adj_325[12]), .n10024(n10024), .n37(n82_adj_325[13]), 
            .n10026(n10026), .n34(n82_adj_325[14]), .n10028(n10028), .\selected_1__N_354[0] (selected_1__N_354[0]), 
            .LM32D_STB_O(LM32D_STB_O), .\LM32I_ADR_O[9] (LM32I_ADR_O[9]), 
            .n41390(n41390), .n30986(n30986), .n47(n47), .\LM32I_ADR_O[14] (LM32I_ADR_O[14]), 
            .\SHAREDBUS_ADR_I[15] (SHAREDBUS_ADR_I[15]), .n41234(n41234), 
            .n61(n61), .bus_error_f_N_1884(bus_error_f_N_1884), .n41429(n41429), 
            .\next_cycle_type[2] (next_cycle_type[2]), .n13990(n13990), 
            .n30900(n30900), .n41410(n41410), .REF_CLK_c_enable_97(REF_CLK_c_enable_97), 
            .\LM32I_ADR_O[11] (LM32I_ADR_O[11]), .n41310(n41310), .n32728(n32728), 
            .\LM32I_ADR_O[13] (LM32I_ADR_O[13]), .ROM_DAT_O({ROM_DAT_O}), 
            .n8(n8_adj_6470), .n8_adj_273(n8_adj_6481), .n8_adj_274(n8_adj_6460), 
            .n8_adj_275(n8_c), .n8_adj_276(n8_adj_6457), .n3(n3_adj_6483), 
            .n3_adj_277(n3_adj_6480), .n8_adj_278(n8_adj_6462), .n3_adj_279(n3_adj_6482), 
            .n8_adj_280(n8_adj_6464), .n8_adj_281(n8_adj_6456), .n3_adj_282(n3_adj_6476), 
            .n8_adj_283(n8_adj_6473), .n8_adj_284(n8_adj_6472), .n8_adj_285(n8_adj_6466), 
            .n8_adj_286(n8_adj_6459), .n8_adj_287(n8_adj_6477), .n3_adj_288(n3_adj_6475), 
            .n41255(n41255), .n15(n15_adj_6526), .n35788(n35788), .n3_adj_289(n3_adj_6474), 
            .n3_adj_290(n3_adj_6471), .n8_adj_291(n8_adj_6469), .n8_adj_292(n8_adj_6468), 
            .n8_adj_293(n8_adj_6467), .n8_adj_294(n8_adj_6465), .LM32D_DAT_O({LM32D_DAT_O}), 
            .n41324(n41324), .data({data}), .n69({n69}), .ebrEBR_DAT_O({ebrEBR_DAT_O}), 
            .\genblk1.write_data_7__N_3573 ({\genblk1.write_data_7__N_3573 }), 
            .n8_adj_296(n8_adj_6463), .n8_adj_297(n8_adj_6461), .n8_adj_298(n8_adj_6458), 
            .n8_adj_299(n8_adj_6455), .n8_adj_300(n8_adj_6454), .n11(n11_adj_6484), 
            .n8_adj_301(n8_adj_6479), .n3_adj_302(n3_adj_6478), .\LM32I_ADR_O[8] (LM32I_ADR_O[8]), 
            .inst3_Empty(inst3_Empty), .n35204(n35204), .\reg_04[29] (reg_04[29]), 
            .n33332(n33332), .\reg_04[4] (reg_04[4]), .n33294(n33294), 
            .\reg_04[14] (reg_04[14]), .n33370(n33370), .\reg_04[17] (reg_04[17]), 
            .n33256(n33256), .\reg_04[22] (reg_04[22]), .n33218(n33218), 
            .\reg_04[24] (reg_04[24]), .n33180(n33180), .n41262(n41262), 
            .n19822(n19822), .\counter[2] (\counter[2] ), .n8_adj_303(n8), 
            .n41344(n41344), .n41345(n41345), .n30231(n30231), .write_enable(write_enable), 
            .\state_1__N_3407[1] (state_1__N_3407[1]), .n6362(n6362), .n41309(n41309), 
            .n87({n87}), .\genblk1.write_data_23__N_3541 ({\genblk1.write_data_23__N_3541 }), 
            .\LM32I_ADR_O[6] (LM32I_ADR_O[6]), .\SHAREDBUS_ADR_I[5] (\SHAREDBUS_ADR_I[5] ), 
            .n41275(n41275), .\LM32I_ADR_O[4] (LM32I_ADR_O[4]), .\SHAREDBUS_ADR_I[29] (\SHAREDBUS_ADR_I[29] ), 
            .n32174(n32174), .\SHAREDBUS_ADR_I[25] (SHAREDBUS_ADR_I[25]), 
            .n35605(n35605), .\SHAREDBUS_ADR_I[20] (SHAREDBUS_ADR_I[20]), 
            .n41289(n41289), .selected({selected_c[1], selected[0]}), 
            .REF_CLK_c(REF_CLK_c), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .\LM32D_ADR_O[10] (LM32D_ADR_O[10]), .n46(n82_adj_325[10]), 
            .n41306(n41306), .\SHAREDBUS_DAT_I[14] (\SHAREDBUS_DAT_I[14] ), 
            .n78({n78}), .\SHAREDBUS_DAT_I[15] (\SHAREDBUS_DAT_I[15] ), 
            .\SHAREDBUS_DAT_I[10] (\SHAREDBUS_DAT_I[10] ), .\SHAREDBUS_DAT_I[9] (\SHAREDBUS_DAT_I[9] ), 
            .\SHAREDBUS_DAT_I[8] (\SHAREDBUS_DAT_I[8] ), .\SHAREDBUS_DAT_I[12] (\SHAREDBUS_DAT_I[12] ), 
            .\SHAREDBUS_DAT_I[11] (\SHAREDBUS_DAT_I[11] ), .n45101(n45101), 
            .\SHAREDBUS_DAT_I[13] (\SHAREDBUS_DAT_I[13] ), .LM32D_CYC_O(LM32D_CYC_O), 
            .n41326(n41326), .locked_N_493(locked_N_493), .REF_CLK_c_enable_1221(REF_CLK_c_enable_1221), 
            .\genblk1.write_data_15__N_3557 ({\genblk1.write_data_15__N_3557 }), 
            .n41292(n41292), .n41488(n41488), .LM32D_SEL_O({LM32D_SEL_O}), 
            .n41307(n41307), .n41485(n41485), .write_ack(write_ack_adj_6523), 
            .n41278(n41278), .n41328(n41328), .\SHAREDBUS_DAT_I[31] (\SHAREDBUS_DAT_I[31] ), 
            .\SHAREDBUS_DAT_I[30] (\SHAREDBUS_DAT_I[30] ), .\SHAREDBUS_DAT_I[24] (\SHAREDBUS_DAT_I[24] ), 
            .\SHAREDBUS_DAT_I[28] (\SHAREDBUS_DAT_I[28] ), .\SHAREDBUS_DAT_I[29] (\SHAREDBUS_DAT_I[29] ), 
            .\LM32D_ADR_O[29] (LM32D_ADR_O[29]), .\LM32I_ADR_O[29] (LM32I_ADR_O[29]), 
            .\LM32D_ADR_O[18] (LM32D_ADR_O[18]), .\LM32I_ADR_O[18] (LM32I_ADR_O[18]), 
            .\SHAREDBUS_ADR_I[18] (SHAREDBUS_ADR_I[18]), .\LM32D_ADR_O[31] (LM32D_ADR_O[31]), 
            .\LM32I_ADR_O[31] (LM32I_ADR_O[31]), .\SHAREDBUS_ADR_I[31] (SHAREDBUS_ADR_I[31]), 
            .\LM32D_ADR_O[27] (LM32D_ADR_O[27]), .\LM32I_ADR_O[27] (LM32I_ADR_O[27]), 
            .\SHAREDBUS_ADR_I[27] (SHAREDBUS_ADR_I[27]), .\LM32D_ADR_O[23] (LM32D_ADR_O[23]), 
            .\LM32I_ADR_O[23] (LM32I_ADR_O[23]), .\SHAREDBUS_ADR_I[23] (\SHAREDBUS_ADR_I[23] ), 
            .\LM32I_ADR_O[10] (LM32I_ADR_O[10]), .\SHAREDBUS_ADR_I[10] (\SHAREDBUS_ADR_I[10] ), 
            .n954({n954}), .\LM32D_ADR_O[15] (LM32D_ADR_O[15]), .\LM32I_ADR_O[15] (LM32I_ADR_O[15]), 
            .\LM32D_ADR_O[26] (LM32D_ADR_O[26]), .\LM32I_ADR_O[26] (LM32I_ADR_O[26]), 
            .\SHAREDBUS_ADR_I[26] (SHAREDBUS_ADR_I[26]), .\LM32D_ADR_O[16] (LM32D_ADR_O[16]), 
            .\LM32I_ADR_O[16] (LM32I_ADR_O[16]), .\SHAREDBUS_ADR_I[16] (SHAREDBUS_ADR_I[16]), 
            .\LM32D_ADR_O[7] (LM32D_ADR_O[7]), .\LM32I_ADR_O[7] (LM32I_ADR_O[7]), 
            .\SHAREDBUS_ADR_I[7] (\SHAREDBUS_ADR_I[7] ), .\LM32D_ADR_O[25] (LM32D_ADR_O[25]), 
            .\LM32I_ADR_O[25] (LM32I_ADR_O[25]), .n953({n953}), .\LM32D_ADR_O[5] (LM32D_ADR_O[5]), 
            .\LM32I_ADR_O[5] (LM32I_ADR_O[5]), .\LM32D_ADR_O[20] (LM32D_ADR_O[20]), 
            .\LM32I_ADR_O[20] (LM32I_ADR_O[20]), .\LM32D_ADR_O[24] (LM32D_ADR_O[24]), 
            .\LM32I_ADR_O[24] (LM32I_ADR_O[24]), .\SHAREDBUS_ADR_I[24] (SHAREDBUS_ADR_I[24]), 
            .\LM32D_ADR_O[22] (LM32D_ADR_O[22]), .\LM32I_ADR_O[22] (LM32I_ADR_O[22]), 
            .\SHAREDBUS_ADR_I[22] (\SHAREDBUS_ADR_I[22] ), .\LM32D_ADR_O[30] (LM32D_ADR_O[30]), 
            .\LM32I_ADR_O[30] (LM32I_ADR_O[30]), .\SHAREDBUS_ADR_I[30] (SHAREDBUS_ADR_I[30]), 
            .\SHAREDBUS_DAT_I[26] (\SHAREDBUS_DAT_I[26] ), .\SHAREDBUS_DAT_I[27] (\SHAREDBUS_DAT_I[27] ), 
            .\SHAREDBUS_DAT_I[25] (\SHAREDBUS_DAT_I[25] ), .write_ack_adj_304(write_ack), 
            .n41243(n41243), .REF_CLK_c_enable_1581(REF_CLK_c_enable_1581), 
            .\LM32D_CTI_O[0] (\LM32D_CTI_O[0] ), .\LM32I_CTI_O[0] (LM32I_CTI_O[0]), 
            .REF_CLK_c_enable_1597(REF_CLK_c_enable_1597), .REF_CLK_c_enable_1605(REF_CLK_c_enable_1605), 
            .REF_CLK_c_enable_1589(REF_CLK_c_enable_1589), .n41329(n41329), 
            .n41387(n41387), .n9(n9_adj_6532), .n12390(n12390), .\LM32D_ADR_O[0] (LM32D_ADR_O[0]), 
            .n71_adj_305(n71), .\LM32D_ADR_O[6] (LM32D_ADR_O[6]), .\LM32D_ADR_O[12] (LM32D_ADR_O[12]), 
            .n41346(n41346), .\LM32I_ADR_O[12] (\LM32I_ADR_O[12] ), .n41303(n41303), 
            .\LM32D_ADR_O[4] (LM32D_ADR_O[4]), .\LM32D_ADR_O[9] (LM32D_ADR_O[9]), 
            .n41347(n41347), .n41222(n41222), .n41304(n41304), .n6034(n6034), 
            .n41330(n41330), .n41331(n41331), .n41332(n41332), .n41333(n41333), 
            .n41334(n41334), .n41335(n41335), .n41336(n41336), .n41337(n41337), 
            .n41338(n41338), .n41339(n41339), .n41193(n41193), .REF_CLK_c_enable_1558(REF_CLK_c_enable_1558), 
            .n41340(n41340), .n41341(n41341), .n41342(n41342), .n41343(n41343), 
            .n96({n96}), .n55(n82_adj_325[7]), .n41279(n41279), .n29830(n29830), 
            .REF_CLK_c_enable_1574(REF_CLK_c_enable_1574), .\genblk1.write_data_31__N_3525 ({\genblk1.write_data_31__N_3525 }), 
            .n41482(n41482), .\LM32I_ADR_O[2] (LM32I_ADR_O[2]), .n32216(n32216), 
            .n61_adj_306(n82_adj_325[5]), .n21(n21_adj_6527), .n33(n33), 
            .n31955(n31955), .n32220(n32220), .n41210(n41210), .n15_adj_307(n15), 
            .n35868(n35868), .n41225(n41225), .n19(n19), .n41226(n41226), 
            .n41260(n41260), .n34816(n34816), .n11831(n11831), .n41323(n41323), 
            .n41239(n41239), .n41238(n41238), .REF_CLK_c_enable_1131(REF_CLK_c_enable_1131), 
            .n41221(n41221), .\LM32D_ADR_O[14] (LM32D_ADR_O[14]), .n41298(n41298), 
            .REF_CLK_c_enable_1550(REF_CLK_c_enable_1550), .REF_CLK_c_enable_1566(REF_CLK_c_enable_1566), 
            .\LM32D_ADR_O[2] (LM32D_ADR_O[2]), .\LM32D_ADR_O[13] (LM32D_ADR_O[13]), 
            .n41300(n41300), .\next_cycle_type[2]_adj_308 (\next_cycle_type[2] ), 
            .\LM32D_ADR_O[11] (LM32D_ADR_O[11]), .n37905(n37905), .n41299(n41299), 
            .n37904(n37904), .\LM32D_ADR_O[8] (LM32D_ADR_O[8]), .n37906(n37906), 
            .n41301(n41301), .n37903(n37903)) /* synthesis syn_module_defined=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(488[1] 529[20])
    lm32_top LM32 (.GND_net(GND_net), .n41300(n41300), .n41194(n41194), 
            .LEDGPIO_ACK_O(LEDGPIO_ACK_O), .n1128(n1096[0]), .REF_CLK_c(REF_CLK_c), 
            .n69({n69}), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .\state_1__N_3407[1] (state_1__N_3407[1]), .ROM_DAT_O({ROM_DAT_O}), 
            .write_enable(write_enable), .n6362(n6362), .n78({n78}), .n87({n87}), 
            .n96({n96}), .\counter[2] (\counter[2] ), .n41246(n41246), 
            .n19808(n19808), .data({data}), .\SHAREDBUS_ADR_I[10] (\SHAREDBUS_ADR_I[10] ), 
            .n41310(n41310), .n41301(n41301), .\SHAREDBUS_ADR_I[7] (\SHAREDBUS_ADR_I[7] ), 
            .n41346(n41346), .\SHAREDBUS_ADR_I[5] (\SHAREDBUS_ADR_I[5] ), 
            .n41347(n41347), .n41344(n41344), .n41345(n41345), .VCC_net(VCC_net), 
            .write_idx_w({write_idx_w}), .n41352(n41352), .n41351(n41351), 
            .w_result({w_result}), .n41350(n41350), .dcache_refill_request(dcache_refill_request), 
            .\operand_1_x[1] (\operand_1_x[1] ), .dc_re(dc_re), .n41430(n41430), 
            .n41432(n41432), .REF_CLK_c_enable_176(REF_CLK_c_enable_176), 
            .n7611(n7611), .n41405(n41405), .REF_CLK_c_enable_164(REF_CLK_c_enable_164), 
            .n41380(n41380), .LM32D_CYC_O(LM32D_CYC_O), .locked_N_493(locked_N_493), 
            .n41356(n41356), .n41355(n41355), .n41353(n41353), .n41358(n41358), 
            .n41359(n41359), .\operand_m[10] (\operand_m[10] ), .\operand_m[9] (\operand_m[9] ), 
            .\operand_m[5] (\operand_m[5] ), .LM32D_WE_O(LM32D_WE_O), .dcache_select_x(dcache_select_x), 
            .n31750(n31750), .n31955(n31955), .n30241(n30241), .n953({n953}), 
            .n41326(n41326), .n41354(n41354), .bie(bie), .n31279(n31279), 
            .\adder_result_x[16] (\adder_result_x[16] ), .\adder_result_x[17] (\adder_result_x[17] ), 
            .\adder_result_x[18] (\adder_result_x[18] ), .\adder_result_x[19] (\adder_result_x[19] ), 
            .\adder_result_x[20] (\adder_result_x[20] ), .\adder_result_x[21] (\adder_result_x[21] ), 
            .\adder_result_x[22] (\adder_result_x[22] ), .\adder_result_x[23] (\adder_result_x[23] ), 
            .\adder_result_x[24] (\adder_result_x[24] ), .\adder_result_x[25] (\adder_result_x[25] ), 
            .\adder_result_x[26] (\adder_result_x[26] ), .\adder_result_x[27] (\adder_result_x[27] ), 
            .\adder_result_x[28] (\adder_result_x[28] ), .\adder_result_x[29] (\adder_result_x[29] ), 
            .\adder_result_x[30] (\adder_result_x[30] ), .\adder_result_x[31] (\adder_result_x[31] ), 
            .n6518(n6518), .n6648(n6648), .bus_error_f_N_1884(bus_error_f_N_1884), 
            .branch_target_d({branch_target_d}), .direction_m(direction_m), 
            .n45103(n45103), .n45099(n45099), .n41394(n41394), .n41401(n41401), 
            .bie_N_3274(bie_N_3274), .pc_f({pc_f}), .n41325(n41325), .n17816(n17816), 
            .n41379(n41379), .\shifter_result_m[21] (\shifter_result_m[21] ), 
            .n41357(n41357), .\left_shift_result[21] (\left_shift_result[21] ), 
            .\left_shift_result[10] (\left_shift_result[10] ), .b({b}), 
            .\p[0] (\p[0] ), .\p[1] (\p[1] ), .\p[2] (\p[2] ), .\p[3] (\p[3] ), 
            .\p[4] (\p[4] ), .\p[5] (\p[5] ), .\p[6] (\p[6] ), .\p[7] (\p[7] ), 
            .\p[8] (\p[8] ), .\p[9] (\p[9] ), .\p[10] (\p[10] ), .\p[11] (\p[11] ), 
            .\p[12] (\p[12] ), .\p[13] (\p[13] ), .\p[14] (\p[14] ), .\p[15] (\p[15] ), 
            .\p[16] (\p[16] ), .\p[17] (\p[17] ), .\p[18] (\p[18] ), .\p[19] (\p[19] ), 
            .\p[20] (\p[20] ), .\p[21] (\p[21] ), .\p[22] (\p[22] ), .\p[23] (\p[23] ), 
            .\p[24] (\p[24] ), .\p[25] (\p[25] ), .\p[26] (\p[26] ), .\p[27] (\p[27] ), 
            .\p[28] (\p[28] ), .\p[29] (\p[29] ), .\p[30] (\p[30] ), .\a[31] (\a[31] ), 
            .t({t}), .LM32D_DAT_O({LM32D_DAT_O}), .REF_CLK_c_enable_1221(REF_CLK_c_enable_1221), 
            .SHAREDBUS_DAT_O({SHAREDBUS_DAT_O}), .LM32D_SEL_O({LM32D_SEL_O}), 
            .\LM32D_ADR_O[0] (LM32D_ADR_O[0]), .\LM32D_CTI_O[0] (\LM32D_CTI_O[0] ), 
            .n38965(n38965), .LM32D_STB_O(LM32D_STB_O), .n21(n21_adj_6527), 
            .\LM32D_ADR_O[1] (LM32D_ADR_O[1]), .\LM32D_ADR_O[2] (LM32D_ADR_O[2]), 
            .\next_cycle_type[2] (\next_cycle_type[2] ), .\LM32D_ADR_O[4] (LM32D_ADR_O[4]), 
            .\LM32D_ADR_O[5] (LM32D_ADR_O[5]), .\d_adr_o_31__N_2278[5] (\d_adr_o_31__N_2278[5] ), 
            .\LM32D_ADR_O[6] (LM32D_ADR_O[6]), .\LM32D_ADR_O[7] (LM32D_ADR_O[7]), 
            .\LM32D_ADR_O[8] (LM32D_ADR_O[8]), .\LM32D_ADR_O[9] (LM32D_ADR_O[9]), 
            .\d_adr_o_31__N_2278[9] (\d_adr_o_31__N_2278[9] ), .\LM32D_ADR_O[10] (LM32D_ADR_O[10]), 
            .\d_adr_o_31__N_2278[10] (\d_adr_o_31__N_2278[10] ), .\LM32D_ADR_O[11] (LM32D_ADR_O[11]), 
            .\LM32D_ADR_O[12] (LM32D_ADR_O[12]), .\LM32D_ADR_O[13] (LM32D_ADR_O[13]), 
            .\LM32D_ADR_O[14] (LM32D_ADR_O[14]), .\LM32D_ADR_O[15] (LM32D_ADR_O[15]), 
            .\LM32D_ADR_O[16] (LM32D_ADR_O[16]), .\LM32D_ADR_O[17] (\LM32D_ADR_O[17] ), 
            .\LM32D_ADR_O[18] (LM32D_ADR_O[18]), .\LM32D_ADR_O[19] (\LM32D_ADR_O[19] ), 
            .\LM32D_ADR_O[20] (LM32D_ADR_O[20]), .\LM32D_ADR_O[21] (LM32D_ADR_O[21]), 
            .\LM32D_ADR_O[22] (LM32D_ADR_O[22]), .\LM32D_ADR_O[23] (LM32D_ADR_O[23]), 
            .\LM32D_ADR_O[24] (LM32D_ADR_O[24]), .\LM32D_ADR_O[25] (LM32D_ADR_O[25]), 
            .\LM32D_ADR_O[26] (LM32D_ADR_O[26]), .\LM32D_ADR_O[27] (LM32D_ADR_O[27]), 
            .\LM32D_ADR_O[28] (LM32D_ADR_O[28]), .\LM32D_ADR_O[29] (LM32D_ADR_O[29]), 
            .\LM32D_ADR_O[30] (LM32D_ADR_O[30]), .\LM32D_ADR_O[31] (LM32D_ADR_O[31]), 
            .n41387(n41387), .n9(n9_adj_6532), .\state[0] (\state[0] ), 
            .\state[2] (\state[2] ), .flush_set({flush_set}), .flush_set_8__N_2513({flush_set_8__N_2513}), 
            .\dcache_refill_address[5] (\dcache_refill_address[5] ), .\dcache_refill_address[9] (\dcache_refill_address[9] ), 
            .\dcache_refill_address[10] (\dcache_refill_address[10] ), .\tmem_write_address[1] (\tmem_write_address[1] ), 
            .\tmem_write_address[5] (\tmem_write_address[5] ), .\tmem_write_address[6] (\tmem_write_address[6] ), 
            .\dmem_write_address[3] (\dmem_write_address[3] ), .\dmem_write_address[7] (\dmem_write_address[7] ), 
            .\dmem_write_address[8] (\dmem_write_address[8] ), .n36337(n36337), 
            .SPI_INT_O_N_4422(SPI_INT_O_N_4422), .SPI_INT_O_N_4417(SPI_INT_O_N_4417), 
            .SPI_INT_O_N_4421(SPI_INT_O_N_4421), .\genblk1.wait_one_tick_done (\genblk1.wait_one_tick_done ), 
            .n6781(n6781), .n6764(n6764), .n6749(n6749), .n41410(n41410), 
            .n13990(n13990), .n32216(n32216), .\LM32I_CTI_O[0] (LM32I_CTI_O[0]), 
            .REF_CLK_c_enable_97(REF_CLK_c_enable_97), .n30900(n30900), 
            .pc_d({pc_d}), .REF_CLK_c_enable_1131(REF_CLK_c_enable_1131), 
            .n6760(n6760), .n45105(n45105), .n73_adj_232(n82_adj_325[1]), 
            .n41461(n41461), .\next_cycle_type[2]_adj_233 (next_cycle_type[2]), 
            .n45080(n45080), .n41390(n41390), .n5223(n5223), .n37955(n37955), 
            .n37956(n37956), .n37954(n37954), .n41250(n41250), .n41251(n41251), 
            .n41279(n41279), .\LM32I_ADR_O[2] (LM32I_ADR_O[2]), .n45079(n45079), 
            .\reg_12[2] (reg_12[2]), .n2(n2_adj_6536), .\reg_12[12] (reg_12[12]), 
            .n40677(n40677), .\reg_12[29] (reg_12[29]), .n2_adj_234(n2_adj_6537), 
            .\reg_12[3] (reg_12[3]), .n2_adj_235(n2_adj_6538), .\reg_12[6] (reg_12[6]), 
            .n2_adj_236(n2_adj_6539), .\reg_12[4] (reg_12[4]), .n2_adj_237(n2_adj_6540), 
            .\reg_12[14] (reg_12[14]), .n2_adj_238(n2_adj_6541), .n41429(n41429), 
            .\reg_12[22] (reg_12[22]), .n2_adj_239(n2_adj_6542), .\reg_12[13] (reg_12[13]), 
            .n2_adj_240(n2_adj_6543), .\reg_12[21] (reg_12[21]), .n2_adj_241(n2_adj_6544), 
            .\reg_12[28] (reg_12[28]), .n2_adj_242(n2_adj_6545), .\reg_12[11] (reg_12[11]), 
            .n2_adj_243(n2_adj_6546), .\reg_12[18] (reg_12[18]), .n2_adj_244(n2_adj_6547), 
            .\reg_12[25] (reg_12[25]), .n2_adj_245(n2_adj_6548), .\reg_12[9] (reg_12[9]), 
            .n2_adj_246(n2_adj_6549), .\reg_12[17] (reg_12[17]), .n2_adj_247(n2_adj_6550), 
            .\reg_12[24] (reg_12[24]), .n2_adj_248(n2_adj_6551), .\reg_12[7] (reg_12[7]), 
            .n2_adj_249(n2_adj_6552), .\reg_12[15] (reg_12[15]), .n2_adj_250(n2_adj_6553), 
            .n6589(n6589), .n6584(n6584), .n37179(n37179), .n6439(n6439), 
            .n6434(n6434), .n37177(n37177), .n6599(n6599), .n6594(n6594), 
            .n37180(n37180), .n6629(n6629), .n6624(n6624), .n37183(n37183), 
            .n6579(n6579), .n6574(n6574), .n37178(n37178), .n6429(n6429), 
            .n6424(n6424), .n37176(n37176), .n6609(n6609), .n6604(n6604), 
            .n37181(n37181), .n6619(n6619), .n6614(n6614), .n37182(n37182), 
            .n37185(n37185), .n37184(n37184), .n37188(n37188), .n37187(n37187), 
            .n37186(n37186), .n37189(n37189), .n7603(n7603), .n7571(n7571), 
            .n7607(n7607), .n7575(n7575), .n7606(n7606), .n7574(n7574), 
            .n7604(n7604), .n7572(n7572), .n7605(n7605), .n7573(n7573), 
            .n7608(n7608), .n7576(n7576), .n7602(n7602), .n7570(n7570), 
            .\selected_1__N_354[0] (selected_1__N_354[0]), .n7601(n7601), 
            .n7569(n7569), .n7600(n7600), .n7568(n7568), .n7599(n7599), 
            .n7567(n7567), .n7598(n7598), .n7566(n7566), .n7597(n7597), 
            .n7565(n7565), .n7596(n7596), .n7564(n7564), .n7595(n7595), 
            .n7563(n7563), .n7594(n7594), .n7562(n7562), .n7593(n7593), 
            .n7561(n7561), .n7592(n7592), .n7560(n7560), .n7584(n7584), 
            .n7552(n7552), .n7583(n7583), .n7551(n7551), .n7582(n7582), 
            .n7550(n7550), .n7581(n7581), .n7549(n7549), .n7580(n7580), 
            .n7548(n7548), .n7579(n7579), .n7547(n7547), .n7578(n7578), 
            .n7546(n7546), .n7577(n7577), .n7545(n7545), .n6750(n6750), 
            .n7591(n7591), .n7559(n7559), .n7590(n7590), .n7558(n7558), 
            .n7589(n7589), .n7557(n7557), .n7588(n7588), .n7556(n7556), 
            .n7587(n7587), .n7555(n7555), .n7586(n7586), .n7554(n7554), 
            .n7585(n7585), .n7553(n7553), .n37501(n37501), .n37500(n37500), 
            .n37502(n37502), .n37499(n37499), .n37498(n37498), .n37497(n37497), 
            .n37496(n37496), .n6751(n6751), .n6752(n6752), .n6753(n6753), 
            .n6754(n6754), .n6755(n6755), .n6756(n6756), .n6757(n6757), 
            .n6758(n6758), .n6759(n6759), .n6761(n6761), .n6762(n6762), 
            .n6763(n6763), .n37495(n37495), .n7672(n7672), .n7640(n7640), 
            .n7673(n7673), .n7641(n7641), .n34(n34_adj_309), .n7674(n7674), 
            .n7642(n7642), .n7675(n7675), .n7643(n7643), .n7676(n7676), 
            .n7644(n7644), .n7671(n7671), .n7639(n7639), .n7670(n7670), 
            .n7638(n7638), .n7669(n7669), .n7637(n7637), .n7668(n7668), 
            .n7636(n7636), .n7667(n7667), .n7635(n7635), .n7666(n7666), 
            .n7634(n7634), .n7665(n7665), .n7633(n7633), .n7664(n7664), 
            .n7632(n7632), .n7663(n7663), .n7631(n7631), .n7662(n7662), 
            .n7630(n7630), .n7661(n7661), .n7629(n7629), .n7660(n7660), 
            .n7628(n7628), .n36(n36), .n7652(n7652), .n7620(n7620), 
            .n7651(n7651), .n7619(n7619), .n7650(n7650), .n7618(n7618), 
            .n7649(n7649), .n7617(n7617), .n37(n37_adj_310), .n7648(n7648), 
            .n7616(n7616), .n7647(n7647), .n7615(n7615), .n7646(n7646), 
            .n7614(n7614), .n7645(n7645), .n7613(n7613), .n7659(n7659), 
            .n7627(n7627), .n7658(n7658), .n7626(n7626), .n7657(n7657), 
            .n7625(n7625), .n7656(n7656), .n7624(n7624), .n7655(n7655), 
            .n7623(n7623), .n7654(n7654), .n7622(n7622), .n7653(n7653), 
            .n7621(n7621), .n37504(n37504), .n37503(n37503), .n37507(n37507), 
            .n37506(n37506), .n37505(n37505), .n37508(n37508), .n45106(n45106), 
            .\LM32I_ADR_O[4] (LM32I_ADR_O[4]), .\LM32I_ADR_O[5] (LM32I_ADR_O[5]), 
            .\LM32I_ADR_O[6] (LM32I_ADR_O[6]), .\LM32I_ADR_O[7] (LM32I_ADR_O[7]), 
            .\LM32I_ADR_O[8] (LM32I_ADR_O[8]), .\LM32I_ADR_O[9] (LM32I_ADR_O[9]), 
            .\LM32I_ADR_O[10] (LM32I_ADR_O[10]), .\LM32I_ADR_O[11] (LM32I_ADR_O[11]), 
            .\LM32I_ADR_O[12] (\LM32I_ADR_O[12] ), .\LM32I_ADR_O[13] (LM32I_ADR_O[13]), 
            .\LM32I_ADR_O[14] (LM32I_ADR_O[14]), .\LM32I_ADR_O[15] (LM32I_ADR_O[15]), 
            .\LM32I_ADR_O[16] (LM32I_ADR_O[16]), .\LM32I_ADR_O[17] (\LM32I_ADR_O[17] ), 
            .\LM32I_ADR_O[18] (LM32I_ADR_O[18]), .\LM32I_ADR_O[19] (\LM32I_ADR_O[19] ), 
            .\LM32I_ADR_O[20] (LM32I_ADR_O[20]), .\LM32I_ADR_O[21] (LM32I_ADR_O[21]), 
            .\LM32I_ADR_O[22] (LM32I_ADR_O[22]), .\LM32I_ADR_O[23] (LM32I_ADR_O[23]), 
            .\LM32I_ADR_O[24] (LM32I_ADR_O[24]), .\LM32I_ADR_O[25] (LM32I_ADR_O[25]), 
            .\LM32I_ADR_O[26] (LM32I_ADR_O[26]), .\LM32I_ADR_O[27] (LM32I_ADR_O[27]), 
            .\LM32I_ADR_O[28] (LM32I_ADR_O[28]), .\LM32I_ADR_O[29] (LM32I_ADR_O[29]), 
            .\LM32I_ADR_O[30] (LM32I_ADR_O[30]), .\LM32I_ADR_O[31] (LM32I_ADR_O[31]), 
            .n949({n949}), .n32220(n32220), .selected({selected_c[1], 
            selected[0]}), .flush_set_adj_272({flush_set_adj_326}), .flush_set_8__N_1953({flush_set_8__N_1953}), 
            .n157({n157}), .n36336(n36336), .n10589(n10589), .n10585(n10585), 
            .n10591(n10591), .n10593(n10593), .n10587(n10587), .n10595(n10595), 
            .n10452(n10452)) /* synthesis syn_module_defined=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(572[2] 613[36])
    \gpio(DATA_WIDTH=32'b01000,INPUT_WIDTH=32'b01,OUTPUT_WIDTH=32'b01,EDGE=1,POSE_EDGE_IRQ=1,INPUT_PORTS_ONLY=0,OUTPUT_PORTS_ONLY=1)  LED (.LEDGPIO_ACK_O(LEDGPIO_ACK_O), 
            .REF_CLK_c(REF_CLK_c), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .PIO_OUT_7__N_3493(PIO_OUT_7__N_3493), .LED_R_c_0(LED_R_c_0), 
            .REF_CLK_c_enable_424(REF_CLK_c_enable_424), .n36338(n36338), 
            .n41345(n41345), .n41344(n41344), .write_ack_N_4033(write_ack_N_4033), 
            .n41185(n41185), .n30156(n30156), .n41347(n41347), .dw10_cs_N_4471(dw10_cs_N_4471), 
            .dw00_cs_N_4467(dw00_cs_N_4467)) /* synthesis syn_module_defined=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(638[2] 654[34])
    \Reg_Comp(reg_08_int_val=32'b010010001101001010101111001101,CLK_MHZ=48.0)  GPO (.LED_G_c_0(LED_G_c_0), 
            .REF_CLK_c(REF_CLK_c), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .n41328(n41328), .\reg_04[0] (reg_04[0]), .write_ack(write_ack), 
            .n35736(n35736), .n15(n15), .n41301(n41301), .n31750(n31750), 
            .n41210(n41210), .n41303(n41303), .n35854(n35854), .n41273(n41273), 
            .n41260(n41260), .n35739(n35739), .n41235(n41235), .\SHAREDBUS_ADR_I[22] (\SHAREDBUS_ADR_I[22] ), 
            .\SHAREDBUS_ADR_I[29] (\SHAREDBUS_ADR_I[29] ), .write_ack_N_4033(write_ack_N_4033), 
            .n41251(n41251), .n41324(n41324), .n41243(n41243), .n41238(n41238), 
            .n41309(n41309), .n41239(n41239), .n41329(n41329), .\GPOout_pins[2] (GPOout_pins[2]), 
            .n41330(n41330), .\GPOout_pins[3] (GPOout_pins[3]), .n41331(n41331), 
            .\GPOout_pins[4] (GPOout_pins[4]), .n41332(n41332), .n41333(n41333), 
            .\GPOout_pins[6] (GPOout_pins[6]), .n41334(n41334), .\GPOout_pins[7] (GPOout_pins[7]), 
            .n41335(n41335), .\SHAREDBUS_DAT_I[8] (\SHAREDBUS_DAT_I[8] ), 
            .\reg_00[9] (reg_00[9]), .\SHAREDBUS_DAT_I[9] (\SHAREDBUS_DAT_I[9] ), 
            .\SHAREDBUS_DAT_I[10] (\SHAREDBUS_DAT_I[10] ), .\reg_00[11] (reg_00[11]), 
            .\SHAREDBUS_DAT_I[11] (\SHAREDBUS_DAT_I[11] ), .\SHAREDBUS_DAT_I[12] (\SHAREDBUS_DAT_I[12] ), 
            .\reg_00[13] (reg_00[13]), .\SHAREDBUS_DAT_I[13] (\SHAREDBUS_DAT_I[13] ), 
            .\reg_00[14] (reg_00[14]), .\SHAREDBUS_DAT_I[14] (\SHAREDBUS_DAT_I[14] ), 
            .\reg_00[15] (reg_00[15]), .\SHAREDBUS_DAT_I[15] (\SHAREDBUS_DAT_I[15] ), 
            .n41336(n41336), .\reg_00[17] (reg_00[17]), .n41337(n41337), 
            .\reg_00[18] (reg_00[18]), .n41338(n41338), .n41339(n41339), 
            .n41340(n41340), .\reg_00[21] (reg_00[21]), .n41341(n41341), 
            .\reg_00[22] (reg_00[22]), .n41342(n41342), .n41343(n41343), 
            .\reg_00[24] (reg_00[24]), .\SHAREDBUS_DAT_I[24] (\SHAREDBUS_DAT_I[24] ), 
            .\reg_00[25] (reg_00[25]), .\SHAREDBUS_DAT_I[25] (\SHAREDBUS_DAT_I[25] ), 
            .\SHAREDBUS_DAT_I[26] (\SHAREDBUS_DAT_I[26] ), .\SHAREDBUS_DAT_I[27] (\SHAREDBUS_DAT_I[27] ), 
            .\reg_00[28] (reg_00[28]), .\SHAREDBUS_DAT_I[28] (\SHAREDBUS_DAT_I[28] ), 
            .\reg_00[29] (reg_00[29]), .\SHAREDBUS_DAT_I[29] (\SHAREDBUS_DAT_I[29] ), 
            .\SHAREDBUS_DAT_I[30] (\SHAREDBUS_DAT_I[30] ), .\SHAREDBUS_DAT_I[31] (\SHAREDBUS_DAT_I[31] ), 
            .n41279(n41279), .n13(n13_adj_6486), .n13_adj_138(n13_adj_6496), 
            .n13_adj_139(n13_adj_6498), .n9(n9_adj_6504), .\reg_04[2] (reg_04[2]), 
            .\reg_04[3] (reg_04[3]), .\reg_04[4] (reg_04[4]), .\reg_04[6] (reg_04[6]), 
            .\reg_04[7] (reg_04[7]), .\reg_04[9] (reg_04[9]), .\reg_04[11] (reg_04[11]), 
            .\reg_04[13] (reg_04[13]), .\reg_04[14] (reg_04[14]), .\reg_04[15] (reg_04[15]), 
            .\reg_04[17] (reg_04[17]), .\reg_04[18] (reg_04[18]), .\reg_04[21] (reg_04[21]), 
            .\reg_04[22] (reg_04[22]), .\reg_04[24] (reg_04[24]), .\reg_04[25] (reg_04[25]), 
            .\reg_04[28] (reg_04[28]), .\reg_04[29] (reg_04[29]), .\GPOwb_DAT_O[8] (GPOwb_DAT_O[8]), 
            .\GPOwb_DAT_O[1] (GPOwb_DAT_O[1]), .n13_adj_140(n13_adj_6490), 
            .n13_adj_141(n13_adj_6492), .n34304(n34304), .n41185(n41185), 
            .n34112(n34112), .\GPOwb_DAT_O[0] (GPOwb_DAT_O[0]), .n11(n11_adj_6494), 
            .n13_adj_142(n13_adj_6500), .\GPOwb_DAT_O[5] (GPOwb_DAT_O[5]), 
            .n13_adj_143(n13_adj_6488), .n13_adj_144(n13_adj_6502), .\SHAREDBUS_ADR_I[20] (SHAREDBUS_ADR_I[20]), 
            .n41242(n41242), .n41250(n41250), .n35577(n35577), .n32366(n32366), 
            .n41310(n41310), .n19(n19), .n41225(n41225), .n35647(n35647), 
            .n41258(n41258), .n35724(n35724), .n41253(n41253), .n41246(n41246), 
            .\SHAREDBUS_ADR_I[26] (SHAREDBUS_ADR_I[26]), .\SHAREDBUS_ADR_I[16] (SHAREDBUS_ADR_I[16]), 
            .n35633(n35633), .read_ack(read_ack), .n41269(n41269), .n34242(n34242), 
            .n41304(n41304), .n33328(n33328), .n33294(n33294), .n32312(n32312), 
            .n33404(n33404), .n33370(n33370), .n33290(n33290), .\SHAREDBUS_ADR_I[24] (SHAREDBUS_ADR_I[24]), 
            .\SHAREDBUS_ADR_I[25] (SHAREDBUS_ADR_I[25]), .\SHAREDBUS_ADR_I[18] (SHAREDBUS_ADR_I[18]), 
            .\SHAREDBUS_ADR_I[27] (SHAREDBUS_ADR_I[27]), .n33256(n33256), 
            .n33252(n33252), .n33218(n33218), .n33214(n33214), .n33180(n33180), 
            .n33356(n33356), .n33366(n33366)) /* synthesis syn_module_defined=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(736[2] 752[34])
    \gpio(DATA_WIDTH=32'b01,INPUT_WIDTH=32'b01,OUTPUT_WIDTH=32'b01,EDGE=1,POSE_EDGE_IRQ=1,INPUT_PORTS_ONLY=0,BOTH_INPUT_AND_OUTPUT=1)  GPIO (.GPIOGPIO_ACK_O(GPIOGPIO_ACK_O), 
            .REF_CLK_c(REF_CLK_c), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .PIO_DATAI_0__N_3822(PIO_DATAI_0__N_3822), .LED_B_c_0(LED_B_c_0), 
            .REF_CLK_c_enable_424(REF_CLK_c_enable_424), .n36339(n36339), 
            .PIO_DATAI({PIO_DATAI}), .n36340(n36340), .n35006(n35006), 
            .PIO_OUT_7__N_3493(PIO_OUT_7__N_3493), .n41275(n41275), .n41310(n41310), 
            .\SHAREDBUS_ADR_I[7] (\SHAREDBUS_ADR_I[7] ), .n954({n954}), 
            .LEDGPIO_ACK_O(LEDGPIO_ACK_O)) /* synthesis syn_module_defined=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(707[2] 724[34])
    \FIFO_Comp(reg_16_int_val=32'b010010001101001010101111001101)  FIFO (.n32828(n32828), 
            .n41246(n41246), .n34372(n34372), .n5223(n5223), .n15(n15), 
            .n41303(n41303), .\SHAREDBUS_ADR_I[25] (SHAREDBUS_ADR_I[25]), 
            .\SHAREDBUS_ADR_I[24] (SHAREDBUS_ADR_I[24]), .\SHAREDBUS_ADR_I[29] (\SHAREDBUS_ADR_I[29] ), 
            .\SHAREDBUS_ADR_I[16] (SHAREDBUS_ADR_I[16]), .n41345(n41345), 
            .\SHAREDBUS_ADR_I[7] (\SHAREDBUS_ADR_I[7] ), .n41186(n41186), 
            .n16(n16_adj_6520), .n17(n17_adj_6393), .n19(n19_adj_6512), 
            .n5(n5_adj_6401), .read_ack(read_ack_adj_6524), .REF_CLK_c(REF_CLK_c), 
            .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), .n31476(n31476), 
            .n19_adj_66(n19_adj_6511), .n5_adj_67(n5), .n16_adj_68(n16_adj_6519), 
            .n17_adj_69(n17_adj_6397), .n16_adj_70(n16_adj_6515), .n22(n22_adj_6405), 
            .n16_adj_71(n16_adj_6514), .n22_adj_72(n22), .n8(n8_adj_6506), 
            .n2(n2_adj_6409), .n16_adj_73(n16_adj_6517), .n22_adj_74(n22_adj_6407), 
            .n16_adj_75(n16_adj_6518), .n22_adj_76(n22_adj_6413), .n8_adj_77(n8_adj_6507), 
            .n2_adj_78(n2_adj_6411), .n41344(n41344), .n19_adj_79(n19_adj_6516), 
            .n26(n26), .n359(n328[1]), .n392(n361[1]), .n16_adj_80(n16_adj_6521), 
            .n17_adj_81(n17_adj_6390), .n16_adj_82(n16_adj_6522), .n17_adj_83(n17_adj_6389), 
            .n17_adj_84(n17_adj_6508), .n5_adj_85(n5_adj_6415), .n13(n13_adj_6453), 
            .n14(n14_adj_6485), .REF_CLK_c_enable_1550(REF_CLK_c_enable_1550), 
            .n41328(n41328), .inst1_FIFOfifo_rst(inst1_FIFOfifo_rst), .REF_CLK_c_enable_1581(REF_CLK_c_enable_1581), 
            .write_ack(write_ack_adj_6523), .write_ack_N_4649(write_ack_N_4649), 
            .inst3_Empty(inst3_Empty), .fiford_reg(fiford_reg), .fiford(fiford), 
            .n40677(n40677), .\SHAREDBUS_ADR_I[23] (\SHAREDBUS_ADR_I[23] ), 
            .\SHAREDBUS_ADR_I[18] (SHAREDBUS_ADR_I[18]), .n32798(n32798), 
            .inst3_Q({inst3_Q}), .n41347(n41347), .n31779(n31779), .n41329(n41329), 
            .n41330(n41330), .n41331(n41331), .n41332(n41332), .n41333(n41333), 
            .n41334(n41334), .n41335(n41335), .REF_CLK_c_enable_1558(REF_CLK_c_enable_1558), 
            .\SHAREDBUS_DAT_I[8] (\SHAREDBUS_DAT_I[8] ), .\SHAREDBUS_DAT_I[9] (\SHAREDBUS_DAT_I[9] ), 
            .\SHAREDBUS_DAT_I[10] (\SHAREDBUS_DAT_I[10] ), .\SHAREDBUS_DAT_I[11] (\SHAREDBUS_DAT_I[11] ), 
            .\SHAREDBUS_DAT_I[12] (\SHAREDBUS_DAT_I[12] ), .\SHAREDBUS_DAT_I[13] (\SHAREDBUS_DAT_I[13] ), 
            .\SHAREDBUS_DAT_I[14] (\SHAREDBUS_DAT_I[14] ), .\SHAREDBUS_DAT_I[15] (\SHAREDBUS_DAT_I[15] ), 
            .REF_CLK_c_enable_1566(REF_CLK_c_enable_1566), .n41336(n41336), 
            .n41337(n41337), .n41338(n41338), .n41339(n41339), .n41340(n41340), 
            .n41341(n41341), .n41342(n41342), .n41343(n41343), .REF_CLK_c_enable_1574(REF_CLK_c_enable_1574), 
            .\SHAREDBUS_DAT_I[24] (\SHAREDBUS_DAT_I[24] ), .\SHAREDBUS_DAT_I[25] (\SHAREDBUS_DAT_I[25] ), 
            .\SHAREDBUS_DAT_I[26] (\SHAREDBUS_DAT_I[26] ), .\SHAREDBUS_DAT_I[27] (\SHAREDBUS_DAT_I[27] ), 
            .\SHAREDBUS_DAT_I[28] (\SHAREDBUS_DAT_I[28] ), .\SHAREDBUS_DAT_I[29] (\SHAREDBUS_DAT_I[29] ), 
            .\SHAREDBUS_DAT_I[30] (\SHAREDBUS_DAT_I[30] ), .\SHAREDBUS_DAT_I[31] (\SHAREDBUS_DAT_I[31] ), 
            .\reg_12[2] (reg_12[2]), .\reg_12[3] (reg_12[3]), .\reg_12[4] (reg_12[4]), 
            .\reg_12[6] (reg_12[6]), .\reg_12[7] (reg_12[7]), .REF_CLK_c_enable_1589(REF_CLK_c_enable_1589), 
            .\reg_12[9] (reg_12[9]), .\reg_12[11] (reg_12[11]), .\reg_12[12] (reg_12[12]), 
            .\reg_12[13] (reg_12[13]), .\reg_12[14] (reg_12[14]), .\reg_12[15] (reg_12[15]), 
            .REF_CLK_c_enable_1597(REF_CLK_c_enable_1597), .\reg_12[17] (reg_12[17]), 
            .\reg_12[18] (reg_12[18]), .\reg_12[21] (reg_12[21]), .\reg_12[22] (reg_12[22]), 
            .\reg_12[24] (reg_12[24]), .REF_CLK_c_enable_1605(REF_CLK_c_enable_1605), 
            .\reg_12[25] (reg_12[25]), .\reg_12[28] (reg_12[28]), .\reg_12[29] (reg_12[29]), 
            .inst3_Full(inst3_Full), .n41193(n41193), .n2_adj_86(n2_adj_6536), 
            .n37903(n37903), .n2_adj_87(n2_adj_6538), .n37905(n37905), 
            .n2_adj_88(n2_adj_6540), .n4893(n4865[4]), .n2_adj_89(n2_adj_6539), 
            .n2_adj_90(n2_adj_6552), .n2_adj_91(n2_adj_6549), .n2_adj_92(n2_adj_6546), 
            .n37904(n37904), .n2_adj_93(n2_adj_6543), .n2_adj_94(n2_adj_6541), 
            .n4883(n4865[14]), .n2_adj_95(n2_adj_6553), .n2_adj_96(n2_adj_6550), 
            .n4880(n4865[17]), .n2_adj_97(n2_adj_6547), .n2_adj_98(n2_adj_6544), 
            .n37906(n37906), .n2_adj_99(n2_adj_6542), .n4875(n4865[22]), 
            .n2_adj_100(n2_adj_6551), .n4873(n4865[24]), .n2_adj_101(n2_adj_6548), 
            .n41275(n41275), .REF_CLK_c_enable_424(REF_CLK_c_enable_424), 
            .n41310(n41310), .n30762(n30762), .n30241(n30241), .n41180(n41180), 
            .n41181(n41181), .\FIFOwb_DAT_O[12] (FIFOwb_DAT_O[12]), .n2_adj_102(n2_adj_6545), 
            .n2_adj_103(n2_adj_6537), .n4868(n4865[29]), .n954({n954}), 
            .n953({n953}), .n41301(n41301), .n32366(n32366), .n41262(n41262), 
            .n41278(n41278), .n35136(n35136), .n33088(n33088), .n41304(n41304), 
            .n34742(n34742), .n41226(n41226), .n41255(n41255), .n41323(n41323), 
            .n5_adj_104(n5_adj_6525), .spiSPI_ACK_O(spiSPI_ACK_O), .n35042(n35042), 
            .n352(n328[8]), .n385(n361[8]), .n19_adj_105(n19_adj_6513), 
            .n26_adj_106(n26_adj_6419), .n19_adj_107(n19_adj_6497), .n25(n25), 
            .n19_adj_108(n19_adj_6505), .n25_adj_109(n25_adj_6433), .n355(n328[5]), 
            .n388(n361[5]), .n19_adj_110(n19_adj_6491), .n5_adj_111(n5_adj_6435), 
            .n19_adj_112(n19_adj_6499), .n25_adj_113(n25_adj_6437), .n17_adj_114(n17_adj_6495), 
            .n22_adj_115(n22_adj_6441), .n8_adj_116(n8_adj_6510), .n2_adj_117(n2_adj_6421), 
            .n19_adj_118(n19_adj_6503), .n25_adj_119(n25_adj_6431), .n19_adj_120(n19_adj_6493), 
            .n25_adj_121(n25_adj_6439), .n360(n328[0]), .n393(n361[0]), 
            .n31183(n31183), .n23(n23), .n31(n31), .n19_adj_122(n19_adj_6489), 
            .n5_adj_123(n5_adj_6428), .n8_adj_124(n8_adj_6509), .n2_adj_125(n2_adj_6417), 
            .n19_adj_126(n19_adj_6501), .n25_adj_127(n25_adj_6443), .n19_adj_128(n19_adj_6487), 
            .n5_adj_129(n5_adj_6424), .n33846(n33846), .\FIFOwb_DAT_O[0] (FIFOwb_DAT_O[0]), 
            .n41210(n41210), .n33864(n33864), .n19_adj_130(n19), .n41258(n41258), 
            .n30949(n30949), .\SHAREDBUS_ADR_I[30] (SHAREDBUS_ADR_I[30]), 
            .n41272(n41272), .n41265(n41265), .n30951(n30951), .n30948(n30948), 
            .n30944(n30944), .\SHAREDBUS_ADR_I[20] (SHAREDBUS_ADR_I[20]), 
            .\SHAREDBUS_ADR_I[26] (SHAREDBUS_ADR_I[26]), .\SHAREDBUS_ADR_I[27] (SHAREDBUS_ADR_I[27]), 
            .\SHAREDBUS_ADR_I[22] (\SHAREDBUS_ADR_I[22] ), .n35844(n35844), 
            .n35866(n35866), .n41274(n41274), .\SHAREDBUS_ADR_I[5] (\SHAREDBUS_ADR_I[5] ), 
            .n41346(n41346), .n41225(n41225), .n35633(n35633), .n35736(n35736), 
            .n41277(n41277), .n41289(n41289), .n32814(n32814), .n35796(n35796), 
            .\FIFOwb_DAT_O[18] (FIFOwb_DAT_O[18]), .\FIFOwb_DAT_O[25] (FIFOwb_DAT_O[25]), 
            .n37954(n37954), .\FIFOwb_DAT_O[31] (FIFOwb_DAT_O[31]), .n37956(n37956), 
            .\FIFOwb_DAT_O[30] (FIFOwb_DAT_O[30]), .n37955(n37955), .\FIFOwb_DAT_O[27] (FIFOwb_DAT_O[27]), 
            .\FIFOwb_DAT_O[26] (FIFOwb_DAT_O[26]), .\FIFOwb_DAT_O[23] (FIFOwb_DAT_O[23]), 
            .\FIFOwb_DAT_O[20] (FIFOwb_DAT_O[20]), .\FIFOwb_DAT_O[19] (FIFOwb_DAT_O[19]), 
            .\FIFOwb_DAT_O[16] (FIFOwb_DAT_O[16]), .\FIFOwb_DAT_O[10] (FIFOwb_DAT_O[10]), 
            .\FIFOwb_DAT_O[8] (FIFOwb_DAT_O[8]), .\FIFOwb_DAT_O[5] (FIFOwb_DAT_O[5]), 
            .\FIFOwb_DAT_O[1] (FIFOwb_DAT_O[1]), .\FIFOwb_DAT_O[21] (FIFOwb_DAT_O[21]), 
            .\FIFOwb_DAT_O[28] (FIFOwb_DAT_O[28]), .\FIFOwb_DAT_O[15] (FIFOwb_DAT_O[15]), 
            .\FIFOwb_DAT_O[13] (FIFOwb_DAT_O[13]), .\FIFOwb_DAT_O[11] (FIFOwb_DAT_O[11]), 
            .\FIFOwb_DAT_O[9] (FIFOwb_DAT_O[9])) /* synthesis syn_module_defined=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(801[2] 824[34])
    
endmodule
//
// Verilog Description of module \spi(SLAVE_NUMBER=32'b01,CLKCNT_WIDTH=16) 
//

module \spi(SLAVE_NUMBER=32'b01,CLKCNT_WIDTH=16)  (sclk_N_5010, IO_SCK_c, 
            spiSPI_ACK_O, REF_CLK_c, REF_CLK_c_enable_1606, spiSPI_DAT_O, 
            rx_shift_data_31__N_4339, n41328, dw10_cs_N_4471, REF_CLK_c_enable_1453, 
            IO_MISO_c, dw00_cs_N_4467, IO_0_c_0, GND_net, VCC_net, 
            IO_MOSI_c, n41329, n41330, n41331, n41332, n41333, n41334, 
            n41335, \SHAREDBUS_DAT_I[8] , \SHAREDBUS_DAT_I[9] , \SHAREDBUS_DAT_I[10] , 
            \SHAREDBUS_DAT_I[11] , \SHAREDBUS_DAT_I[12] , \SHAREDBUS_DAT_I[13] , 
            \SHAREDBUS_DAT_I[14] , \SHAREDBUS_DAT_I[15] , n41336, n41337, 
            n41338, n41339, n41340, n41341, n41342, n41343, \SHAREDBUS_DAT_I[24] , 
            \SHAREDBUS_DAT_I[25] , \SHAREDBUS_DAT_I[26] , \SHAREDBUS_DAT_I[27] , 
            \SHAREDBUS_DAT_I[28] , \SHAREDBUS_DAT_I[29] , \SHAREDBUS_DAT_I[30] , 
            \SHAREDBUS_DAT_I[31] , n45179, n41225, \LM32D_ADR_O[1] , 
            n41380, \LM32D_ADR_O[0] , n30156, n41246, n30986, n41310, 
            n41304, n35042, \inst_reg[15] , n10865, n41191, n41345, 
            n41344, n41347, n34742, SPI_INT_O_N_4422, SPI_INT_O_N_4417, 
            SPI_INT_O_N_4421, n953, n954, n34304, \genblk1.wait_one_tick_done ) /* synthesis syn_module_defined=1 */ ;
    output sclk_N_5010;
    output IO_SCK_c;
    output spiSPI_ACK_O;
    input REF_CLK_c;
    input REF_CLK_c_enable_1606;
    output [31:0]spiSPI_DAT_O;
    output rx_shift_data_31__N_4339;
    input n41328;
    input dw10_cs_N_4471;
    output REF_CLK_c_enable_1453;
    input IO_MISO_c;
    input dw00_cs_N_4467;
    output IO_0_c_0;
    input GND_net;
    input VCC_net;
    output IO_MOSI_c;
    input n41329;
    input n41330;
    input n41331;
    input n41332;
    input n41333;
    input n41334;
    input n41335;
    input \SHAREDBUS_DAT_I[8] ;
    input \SHAREDBUS_DAT_I[9] ;
    input \SHAREDBUS_DAT_I[10] ;
    input \SHAREDBUS_DAT_I[11] ;
    input \SHAREDBUS_DAT_I[12] ;
    input \SHAREDBUS_DAT_I[13] ;
    input \SHAREDBUS_DAT_I[14] ;
    input \SHAREDBUS_DAT_I[15] ;
    input n41336;
    input n41337;
    input n41338;
    input n41339;
    input n41340;
    input n41341;
    input n41342;
    input n41343;
    input \SHAREDBUS_DAT_I[24] ;
    input \SHAREDBUS_DAT_I[25] ;
    input \SHAREDBUS_DAT_I[26] ;
    input \SHAREDBUS_DAT_I[27] ;
    input \SHAREDBUS_DAT_I[28] ;
    input \SHAREDBUS_DAT_I[29] ;
    input \SHAREDBUS_DAT_I[30] ;
    input \SHAREDBUS_DAT_I[31] ;
    output n45179;
    input n41225;
    input \LM32D_ADR_O[1] ;
    input n41380;
    input \LM32D_ADR_O[0] ;
    output n30156;
    input n41246;
    input n30986;
    input n41310;
    input n41304;
    input n35042;
    input \inst_reg[15] ;
    input n10865;
    output n41191;
    input n41345;
    input n41344;
    input n41347;
    input n34742;
    output SPI_INT_O_N_4422;
    output SPI_INT_O_N_4417;
    output SPI_INT_O_N_4421;
    input [0:0]n953;
    input [0:0]n954;
    output n34304;
    input \genblk1.wait_one_tick_done ;
    
    wire sclk_N_5010 /* synthesis is_inv_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(57[11:19])
    wire IO_SCK_c /* synthesis is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(28[3:9])
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    
    wire n31773, reg_rd;
    wire [31:0]SPI_DAT_O_31__N_4307;
    wire [31:0]reg_rxdata;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(148[28:38])
    
    wire rx_latch_flag;
    wire [31:0]rx_shift_data;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(150[28:41])
    wire [31:0]reg_txdata;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(149[28:38])
    
    wire reg_txdata_31__N_4306;
    wire [31:0]latch_s_data;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(147[28:40])
    wire [2:0]\genblk1.c_status ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(269[28:36])
    
    wire n41383, n11367;
    wire [5:0]\genblk1.data_cnt ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(267[28:36])
    
    wire n10, n41423;
    wire [15:0]n69;
    wire [15:0]n87;
    
    wire dw04_cs, dw04_cs_N_4468, dw08_cs, dw08_cs_N_4469, dw0c_cs, 
        dw0c_cs_N_4470, dw10_cs, reg_wr, reg_wr_N_4472, reg_rd_N_4474;
    wire [2:0]\genblk1.n_status_2__N_4368 ;
    
    wire n12376;
    wire [2:0]\genblk1.n_status ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(270[28:36])
    
    wire SCLK_MASTER_N_4428, rx_latch_flag_N_4481;
    wire [8:0]reg_status;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(162[28:38])
    
    wire n12374, REF_CLK_c_enable_73, reg_status_4__N_4268, n12382, 
        REF_CLK_c_enable_74, reg_status_7__N_4251, reg_status_5__N_4266, 
        dw00_cs, SS_N_4105, n12, REF_CLK_c_enable_1229, n15969, n41297, 
        n11393, n6264, read_wait_done, n6364, n27517;
    wire [15:0]\genblk1.clock_cnt ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(266[28:37])
    
    wire n27516, n31905, n31971, n12_adj_6337;
    wire [10:0]reg_control;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(154[28:39])
    
    wire reg_control_10__N_4245, REF_CLK_c_enable_760, n9228, n17939, 
        n3, n36490;
    wire [0:0]\genblk1.reg_ssmask ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(265[28:38])
    
    wire \genblk1.reg_ssmask_0__N_4110 , n38969, n27515, n38970, n27514;
    wire [7:0]n4962;
    wire [31:0]n324;
    
    wire n27513, n27512, n27511, n27510;
    wire [31:0]tx_shift_data;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(151[28:41])
    wire [31:0]tx_shift_data_31__N_4212;
    
    wire n35090, n12424, n12422, n28997, n12418, n9, n35244;
    wire [2:0]\genblk1.n_status_2__N_4362 ;
    
    wire n29807, n9215, n1, n35472, n7707, n41442, rx_latch_flag_N_4482;
    wire [2:0]\genblk1.n_status_2__N_4302 ;
    
    wire \genblk1.n_status_2__N_4305 , n3_adj_6338, n6, n35350, n35246, 
        reg_status_6__N_4260, reg_status_7__N_4253, n12_adj_6339, n41209, 
        n1_adj_6340, n35456, n41406, n35254, SPI_INT_O_N_4420, n35354, 
        n6019, n5, n35468, n41422, n34628, n34618, n34620, n34606, 
        n34610, n34604;
    
    INV i35876 (.A(IO_SCK_c), .Z(sclk_N_5010));
    FD1S3DX SPI_ACK_O_254 (.D(n31773), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(spiSPI_ACK_O)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(247[10] 250[25])
    defparam SPI_ACK_O_254.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i0 (.D(SPI_DAT_O_31__N_4307[0]), .SP(reg_rd), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i0.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i0 (.D(rx_shift_data[0]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i0.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i0 (.D(latch_s_data[0]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i0.GSR = "ENABLED";
    LUT4 i33280_3_lut_4_lut (.A(\genblk1.c_status [1]), .B(n41383), .C(IO_SCK_c), 
         .D(n11367), .Z(rx_shift_data_31__N_4339)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(431[17:38])
    defparam i33280_3_lut_4_lut.init = 16'h0002;
    FD1S3DX \genblk1.data_cnt__i0  (.D(n10), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.data_cnt [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(402[12] 411[35])
    defparam \genblk1.data_cnt__i0 .GSR = "ENABLED";
    LUT4 i14803_2_lut_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(n41423), 
         .C(n69[0]), .D(n11367), .Z(n87[0])) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i14803_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i15254_2_lut_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(n41423), 
         .C(n69[1]), .D(n11367), .Z(n87[1])) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i15254_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i15255_2_lut_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(n41423), 
         .C(n69[2]), .D(n11367), .Z(n87[2])) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i15255_2_lut_3_lut_4_lut.init = 16'he000;
    FD1S3DX latch_s_data_i0 (.D(n41328), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i0.GSR = "ENABLED";
    FD1S3DX dw04_cs_239 (.D(dw04_cs_N_4468), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(dw04_cs)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(180[15] 186[9])
    defparam dw04_cs_239.GSR = "ENABLED";
    FD1S3DX dw08_cs_240 (.D(dw08_cs_N_4469), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(dw08_cs)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(180[15] 186[9])
    defparam dw08_cs_240.GSR = "ENABLED";
    FD1S3DX dw0c_cs_241 (.D(dw0c_cs_N_4470), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(dw0c_cs)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(180[15] 186[9])
    defparam dw0c_cs_241.GSR = "ENABLED";
    FD1S3DX dw10_cs_242 (.D(dw10_cs_N_4471), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(dw10_cs)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(180[15] 186[9])
    defparam dw10_cs_242.GSR = "ENABLED";
    FD1S3DX reg_wr_243 (.D(reg_wr_N_4472), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(reg_wr)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(192[15] 195[9])
    defparam reg_wr_243.GSR = "ENABLED";
    FD1S3DX reg_rd_244 (.D(reg_rd_N_4474), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(reg_rd)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(192[15] 195[9])
    defparam reg_rd_244.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i0 (.D(IO_MISO_c), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i0.GSR = "ENABLED";
    FD1S3DX \genblk1.pending_data_256  (.D(n12376), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.n_status_2__N_4368 [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(277[11] 280[49])
    defparam \genblk1.pending_data_256 .GSR = "ENABLED";
    FD1S3DX \genblk1.c_status_i0  (.D(\genblk1.n_status [0]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.c_status [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(349[10:31])
    defparam \genblk1.c_status_i0 .GSR = "ENABLED";
    FD1S3DX SCLK_MASTER_261 (.D(SCLK_MASTER_N_4428), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(IO_SCK_c)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(314[11] 315[46])
    defparam SCLK_MASTER_261.GSR = "ENABLED";
    LUT4 i15256_2_lut_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(n41423), 
         .C(n69[3]), .D(n11367), .Z(n87[3])) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i15256_2_lut_3_lut_4_lut.init = 16'he000;
    FD1S3DX rx_latch_flag_263 (.D(rx_latch_flag_N_4481), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(rx_latch_flag)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(331[12] 334[32])
    defparam rx_latch_flag_263.GSR = "ENABLED";
    FD1S3BX reg_trdy_273 (.D(n12374), .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), 
            .Q(reg_status[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(449[12] 452[24])
    defparam reg_trdy_273.GSR = "ENABLED";
    FD1P3DX reg_toe_274 (.D(reg_status_4__N_4268), .SP(REF_CLK_c_enable_73), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_status[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(457[12] 460[26])
    defparam reg_toe_274.GSR = "ENABLED";
    FD1S3DX reg_rrdy_275 (.D(n12382), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(reg_status[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(466[12] 475[31])
    defparam reg_rrdy_275.GSR = "ENABLED";
    FD1P3DX reg_roe_276 (.D(reg_status_7__N_4251), .SP(REF_CLK_c_enable_74), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_status[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(466[12] 475[31])
    defparam reg_roe_276.GSR = "ENABLED";
    FD1S3BX reg_tmt_277 (.D(reg_status_5__N_4266), .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), 
            .Q(reg_status[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(480[12] 483[26])
    defparam reg_tmt_277.GSR = "ENABLED";
    FD1S3DX dw00_cs_238 (.D(dw00_cs_N_4467), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(dw00_cs)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(180[15] 186[9])
    defparam dw00_cs_238.GSR = "ENABLED";
    FD1S3BX SS_N_MASTER_0__260 (.D(SS_N_4105), .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), 
            .Q(IO_0_c_0)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(302[11] 307[45])
    defparam SS_N_MASTER_0__260.GSR = "ENABLED";
    LUT4 i15257_2_lut_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(n41423), 
         .C(n69[4]), .D(n11367), .Z(n87[4])) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i15257_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i15258_2_lut_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(n41423), 
         .C(n69[5]), .D(n11367), .Z(n87[5])) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i15258_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i15259_2_lut_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(n41423), 
         .C(n69[6]), .D(n11367), .Z(n87[6])) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i15259_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i15260_2_lut_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(n41423), 
         .C(n69[7]), .D(n11367), .Z(n87[7])) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i15260_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i15261_2_lut_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(n41423), 
         .C(n69[8]), .D(n11367), .Z(n87[8])) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i15261_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i15262_2_lut_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(n41423), 
         .C(n69[9]), .D(n11367), .Z(n87[9])) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i15262_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i15263_2_lut_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(n41423), 
         .C(n69[10]), .D(n11367), .Z(n87[10])) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i15263_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i15264_2_lut_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(n41423), 
         .C(n69[11]), .D(n11367), .Z(n87[11])) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i15264_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i15265_2_lut_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(n41423), 
         .C(n69[12]), .D(n11367), .Z(n87[12])) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i15265_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i15266_2_lut_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(n41423), 
         .C(n69[13]), .D(n11367), .Z(n87[13])) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i15266_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i15267_2_lut_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(n41423), 
         .C(n69[14]), .D(n11367), .Z(n87[14])) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i15267_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i15525_2_lut_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(n41423), 
         .C(n69[15]), .D(n11367), .Z(n87[15])) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i15525_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i1_2_lut_rep_818 (.A(n11367), .B(n12), .Z(REF_CLK_c_enable_1229)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_rep_818.init = 16'h4444;
    LUT4 i24_3_lut_4_lut (.A(n11367), .B(n12), .C(n15969), .D(\genblk1.data_cnt [0]), 
         .Z(n10)) /* synthesis lut_function=(A (D)+!A !(B (C+(D))+!B !(D))) */ ;
    defparam i24_3_lut_4_lut.init = 16'hbb04;
    LUT4 i1_3_lut_4_lut (.A(n11367), .B(n41297), .C(n11393), .D(n15969), 
         .Z(n6264)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[16:38])
    defparam i1_3_lut_4_lut.init = 16'hff10;
    FD1S3DX read_wait_done_255 (.D(n6364), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(read_wait_done)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(256[10] 259[30])
    defparam read_wait_done_255.GSR = "ENABLED";
    LUT4 mux_70_i32_4_lut (.A(reg_txdata[31]), .B(reg_rxdata[31]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i32_4_lut.init = 16'hcac0;
    LUT4 mux_70_i31_4_lut (.A(reg_txdata[30]), .B(reg_rxdata[30]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i31_4_lut.init = 16'hcac0;
    FD1P3DX reg_rxdata_i0_i31 (.D(rx_shift_data[31]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i31.GSR = "ENABLED";
    LUT4 mux_70_i30_4_lut (.A(reg_txdata[29]), .B(reg_rxdata[29]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i30_4_lut.init = 16'hcac0;
    FD1P3DX reg_rxdata_i0_i30 (.D(rx_shift_data[30]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i30.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i29 (.D(rx_shift_data[29]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i29.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i28 (.D(rx_shift_data[28]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i28.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i27 (.D(rx_shift_data[27]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i27.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i26 (.D(rx_shift_data[26]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i26.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i25 (.D(rx_shift_data[25]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i25.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i24 (.D(rx_shift_data[24]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i24.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i23 (.D(rx_shift_data[23]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i23.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i22 (.D(rx_shift_data[22]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i22.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i21 (.D(rx_shift_data[21]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i21.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i20 (.D(rx_shift_data[20]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i20.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i19 (.D(rx_shift_data[19]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i19.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i18 (.D(rx_shift_data[18]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i18.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i17 (.D(rx_shift_data[17]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i17.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i16 (.D(rx_shift_data[16]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i16.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i15 (.D(rx_shift_data[15]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i15.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i14 (.D(rx_shift_data[14]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i14.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i13 (.D(rx_shift_data[13]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i13.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i12 (.D(rx_shift_data[12]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i12.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i11 (.D(rx_shift_data[11]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i11.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i10 (.D(rx_shift_data[10]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i10.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i9 (.D(rx_shift_data[9]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i9.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i8 (.D(rx_shift_data[8]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i8.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i7 (.D(rx_shift_data[7]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i7.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i6 (.D(rx_shift_data[6]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i6.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i5 (.D(rx_shift_data[5]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i5.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i4 (.D(rx_shift_data[4]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i4.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i3 (.D(rx_shift_data[3]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i3.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i2 (.D(rx_shift_data[2]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i2.GSR = "ENABLED";
    FD1P3DX reg_rxdata_i0_i1 (.D(rx_shift_data[1]), .SP(rx_latch_flag), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_rxdata[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(207[11] 208[53])
    defparam reg_rxdata_i0_i1.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i31 (.D(SPI_DAT_O_31__N_4307[31]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i31.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i30 (.D(SPI_DAT_O_31__N_4307[30]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i30.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i29 (.D(SPI_DAT_O_31__N_4307[29]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i29.GSR = "ENABLED";
    LUT4 mux_70_i29_4_lut (.A(reg_txdata[28]), .B(reg_rxdata[28]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[28])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i29_4_lut.init = 16'hcac0;
    FD1P3DX SPI_DAT_O_i0_i28 (.D(SPI_DAT_O_31__N_4307[28]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i28.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i27 (.D(SPI_DAT_O_31__N_4307[27]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i27.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i26 (.D(SPI_DAT_O_31__N_4307[26]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i26.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i25 (.D(SPI_DAT_O_31__N_4307[25]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i25.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i24 (.D(SPI_DAT_O_31__N_4307[24]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i24.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i23 (.D(SPI_DAT_O_31__N_4307[23]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i23.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i22 (.D(SPI_DAT_O_31__N_4307[22]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i22.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i21 (.D(SPI_DAT_O_31__N_4307[21]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i21.GSR = "ENABLED";
    LUT4 mux_70_i28_4_lut (.A(reg_txdata[27]), .B(reg_rxdata[27]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[27])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i28_4_lut.init = 16'hcac0;
    FD1P3DX SPI_DAT_O_i0_i20 (.D(SPI_DAT_O_31__N_4307[20]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i20.GSR = "ENABLED";
    LUT4 mux_70_i27_4_lut (.A(reg_txdata[26]), .B(reg_rxdata[26]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[26])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i27_4_lut.init = 16'hcac0;
    FD1P3DX SPI_DAT_O_i0_i19 (.D(SPI_DAT_O_31__N_4307[19]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i19.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i18 (.D(SPI_DAT_O_31__N_4307[18]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i18.GSR = "ENABLED";
    LUT4 mux_70_i26_4_lut (.A(reg_txdata[25]), .B(reg_rxdata[25]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[25])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i26_4_lut.init = 16'hcac0;
    LUT4 mux_70_i25_4_lut (.A(reg_txdata[24]), .B(reg_rxdata[24]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[24])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i25_4_lut.init = 16'hcac0;
    LUT4 mux_70_i24_4_lut (.A(reg_txdata[23]), .B(reg_rxdata[23]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i24_4_lut.init = 16'hcac0;
    FD1P3DX SPI_DAT_O_i0_i17 (.D(SPI_DAT_O_31__N_4307[17]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i17.GSR = "ENABLED";
    CCU2C \genblk1.clock_cnt_2249_add_4_17  (.A0(\genblk1.clock_cnt [15]), 
          .B0(GND_net), .C0(GND_net), .D0(VCC_net), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27517), .S0(n69[15]));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249_add_4_17 .INIT0 = 16'haaa0;
    defparam \genblk1.clock_cnt_2249_add_4_17 .INIT1 = 16'h0000;
    defparam \genblk1.clock_cnt_2249_add_4_17 .INJECT1_0 = "NO";
    defparam \genblk1.clock_cnt_2249_add_4_17 .INJECT1_1 = "NO";
    LUT4 mux_70_i23_4_lut (.A(reg_txdata[22]), .B(reg_rxdata[22]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i23_4_lut.init = 16'hcac0;
    CCU2C \genblk1.clock_cnt_2249_add_4_15  (.A0(\genblk1.clock_cnt [13]), 
          .B0(GND_net), .C0(GND_net), .D0(VCC_net), .A1(\genblk1.clock_cnt [14]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n27516), .COUT(n27517), 
          .S0(n69[13]), .S1(n69[14]));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249_add_4_15 .INIT0 = 16'haaa0;
    defparam \genblk1.clock_cnt_2249_add_4_15 .INIT1 = 16'haaa0;
    defparam \genblk1.clock_cnt_2249_add_4_15 .INJECT1_0 = "NO";
    defparam \genblk1.clock_cnt_2249_add_4_15 .INJECT1_1 = "NO";
    PFUMX i23 (.BLUT(n31905), .ALUT(n31971), .C0(\genblk1.data_cnt [1]), 
          .Z(n12_adj_6337));
    LUT4 mux_70_i22_4_lut (.A(reg_txdata[21]), .B(reg_rxdata[21]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i22_4_lut.init = 16'hcac0;
    FD1P3DX reg_ie_252 (.D(latch_s_data[8]), .SP(reg_control_10__N_4245), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_control[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(230[10] 236[50])
    defparam reg_ie_252.GSR = "ENABLED";
    FD1P3DX reg_sso_253 (.D(latch_s_data[10]), .SP(reg_control_10__N_4245), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_control[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(230[10] 236[50])
    defparam reg_sso_253.GSR = "ENABLED";
    FD1P3DX MOSI_MASTER_271 (.D(n9228), .SP(REF_CLK_c_enable_760), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(IO_MOSI_c)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam MOSI_MASTER_271.GSR = "ENABLED";
    FD1P3DX reg_itrdy_250 (.D(latch_s_data[6]), .SP(reg_control_10__N_4245), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_control[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(230[10] 236[50])
    defparam reg_itrdy_250.GSR = "ENABLED";
    PFUMX i8 (.BLUT(n17939), .ALUT(n3), .C0(n36490), .Z(SPI_DAT_O_31__N_4307[8]));
    FD1P3DX reg_iroe_248 (.D(latch_s_data[3]), .SP(reg_control_10__N_4245), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_control[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(230[10] 236[50])
    defparam reg_iroe_248.GSR = "ENABLED";
    FD1P3DX reg_itoe_249 (.D(latch_s_data[4]), .SP(reg_control_10__N_4245), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_control[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(230[10] 236[50])
    defparam reg_itoe_249.GSR = "ENABLED";
    FD1P3DX \genblk1.reg_ssmask_0__258  (.D(latch_s_data[0]), .SP(\genblk1.reg_ssmask_0__N_4110 ), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\genblk1.reg_ssmask [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(296[11] 297[62])
    defparam \genblk1.reg_ssmask_0__258 .GSR = "ENABLED";
    FD1P3DX reg_irrdy_251 (.D(latch_s_data[7]), .SP(reg_control_10__N_4245), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_control[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(230[10] 236[50])
    defparam reg_irrdy_251.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i16 (.D(SPI_DAT_O_31__N_4307[16]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i16.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i15 (.D(SPI_DAT_O_31__N_4307[15]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i15.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i14 (.D(SPI_DAT_O_31__N_4307[14]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i14.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i13 (.D(SPI_DAT_O_31__N_4307[13]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i13.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i12 (.D(SPI_DAT_O_31__N_4307[12]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i12.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i11 (.D(SPI_DAT_O_31__N_4307[11]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i11.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i10 (.D(SPI_DAT_O_31__N_4307[10]), .SP(reg_rd), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i10.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i9 (.D(SPI_DAT_O_31__N_4307[9]), .SP(reg_rd), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i9.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i8 (.D(SPI_DAT_O_31__N_4307[8]), .SP(reg_rd), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i8.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i7 (.D(SPI_DAT_O_31__N_4307[7]), .SP(reg_rd), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i7.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i6 (.D(SPI_DAT_O_31__N_4307[6]), .SP(reg_rd), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i6.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i5 (.D(SPI_DAT_O_31__N_4307[5]), .SP(reg_rd), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i5.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i4 (.D(SPI_DAT_O_31__N_4307[4]), .SP(reg_rd), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i4.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i3 (.D(SPI_DAT_O_31__N_4307[3]), .SP(reg_rd), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i3.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i2 (.D(SPI_DAT_O_31__N_4307[2]), .SP(reg_rd), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i2.GSR = "ENABLED";
    FD1P3DX SPI_DAT_O_i0_i1 (.D(SPI_DAT_O_31__N_4307[1]), .SP(reg_rd), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(spiSPI_DAT_O[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(285[11] 291[48])
    defparam SPI_DAT_O_i0_i1.GSR = "ENABLED";
    LUT4 \genblk1.n_status_1__bdd_4_lut_33567  (.A(\genblk1.n_status [1]), 
         .B(\genblk1.c_status [1]), .C(\genblk1.c_status [0]), .D(n11367), 
         .Z(n38969)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam \genblk1.n_status_1__bdd_4_lut_33567 .init = 16'h0200;
    CCU2C \genblk1.clock_cnt_2249_add_4_13  (.A0(\genblk1.clock_cnt [11]), 
          .B0(GND_net), .C0(GND_net), .D0(VCC_net), .A1(\genblk1.clock_cnt [12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n27515), .COUT(n27516), 
          .S0(n69[11]), .S1(n69[12]));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249_add_4_13 .INIT0 = 16'haaa0;
    defparam \genblk1.clock_cnt_2249_add_4_13 .INIT1 = 16'haaa0;
    defparam \genblk1.clock_cnt_2249_add_4_13 .INJECT1_0 = "NO";
    defparam \genblk1.clock_cnt_2249_add_4_13 .INJECT1_1 = "NO";
    LUT4 \genblk1.n_status_1__bdd_4_lut  (.A(n11393), .B(\genblk1.c_status [1]), 
         .C(\genblk1.c_status [0]), .D(n11367), .Z(n38970)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C))+!A (B+(C))) */ ;
    defparam \genblk1.n_status_1__bdd_4_lut .init = 16'hfc7c;
    FD1S3DX \genblk1.clock_cnt_2249__i0  (.D(n87[0]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.clock_cnt [0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249__i0 .GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i1 (.D(latch_s_data[1]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i1.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i2 (.D(latch_s_data[2]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i2.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i3 (.D(latch_s_data[3]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i3.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i4 (.D(latch_s_data[4]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i4.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i5 (.D(latch_s_data[5]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i5.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i6 (.D(latch_s_data[6]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i6.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i7 (.D(latch_s_data[7]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i7.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i8 (.D(latch_s_data[8]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i8.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i9 (.D(latch_s_data[9]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i9.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i10 (.D(latch_s_data[10]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i10.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i11 (.D(latch_s_data[11]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i11.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i12 (.D(latch_s_data[12]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i12.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i13 (.D(latch_s_data[13]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i13.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i14 (.D(latch_s_data[14]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i14.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i15 (.D(latch_s_data[15]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i15.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i16 (.D(latch_s_data[16]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i16.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i17 (.D(latch_s_data[17]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i17.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i18 (.D(latch_s_data[18]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i18.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i19 (.D(latch_s_data[19]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i19.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i20 (.D(latch_s_data[20]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i20.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i21 (.D(latch_s_data[21]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i21.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i22 (.D(latch_s_data[22]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i22.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i23 (.D(latch_s_data[23]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i23.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i24 (.D(latch_s_data[24]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i24.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i25 (.D(latch_s_data[25]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i25.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i26 (.D(latch_s_data[26]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i26.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i27 (.D(latch_s_data[27]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i27.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i28 (.D(latch_s_data[28]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i28.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i29 (.D(latch_s_data[29]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i29.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i30 (.D(latch_s_data[30]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i30.GSR = "ENABLED";
    FD1P3DX reg_txdata_i0_i31 (.D(latch_s_data[31]), .SP(reg_txdata_31__N_4306), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_txdata[31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[11] 215[55])
    defparam reg_txdata_i0_i31.GSR = "ENABLED";
    CCU2C \genblk1.clock_cnt_2249_add_4_11  (.A0(\genblk1.clock_cnt [9]), 
          .B0(GND_net), .C0(GND_net), .D0(VCC_net), .A1(\genblk1.clock_cnt [10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n27514), .COUT(n27515), 
          .S0(n69[9]), .S1(n69[10]));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249_add_4_11 .INIT0 = 16'haaa0;
    defparam \genblk1.clock_cnt_2249_add_4_11 .INIT1 = 16'haaa0;
    defparam \genblk1.clock_cnt_2249_add_4_11 .INJECT1_0 = "NO";
    defparam \genblk1.clock_cnt_2249_add_4_11 .INJECT1_1 = "NO";
    PFUMX mux_70_i8 (.BLUT(n4962[5]), .ALUT(n324[7]), .C0(n36490), .Z(SPI_DAT_O_31__N_4307[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;
    CCU2C \genblk1.clock_cnt_2249_add_4_9  (.A0(\genblk1.clock_cnt [7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\genblk1.clock_cnt [8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n27513), .COUT(n27514), .S0(n69[7]), 
          .S1(n69[8]));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249_add_4_9 .INIT0 = 16'haaa0;
    defparam \genblk1.clock_cnt_2249_add_4_9 .INIT1 = 16'haaa0;
    defparam \genblk1.clock_cnt_2249_add_4_9 .INJECT1_0 = "NO";
    defparam \genblk1.clock_cnt_2249_add_4_9 .INJECT1_1 = "NO";
    PFUMX mux_70_i7 (.BLUT(n4962[4]), .ALUT(n324[6]), .C0(n36490), .Z(SPI_DAT_O_31__N_4307[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;
    CCU2C \genblk1.clock_cnt_2249_add_4_7  (.A0(\genblk1.clock_cnt [5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\genblk1.clock_cnt [6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n27512), .COUT(n27513), .S0(n69[5]), 
          .S1(n69[6]));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249_add_4_7 .INIT0 = 16'haaa0;
    defparam \genblk1.clock_cnt_2249_add_4_7 .INIT1 = 16'haaa0;
    defparam \genblk1.clock_cnt_2249_add_4_7 .INJECT1_0 = "NO";
    defparam \genblk1.clock_cnt_2249_add_4_7 .INJECT1_1 = "NO";
    CCU2C \genblk1.clock_cnt_2249_add_4_5  (.A0(\genblk1.clock_cnt [3]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\genblk1.clock_cnt [4]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n27511), .COUT(n27512), .S0(n69[3]), 
          .S1(n69[4]));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249_add_4_5 .INIT0 = 16'haaa0;
    defparam \genblk1.clock_cnt_2249_add_4_5 .INIT1 = 16'haaa0;
    defparam \genblk1.clock_cnt_2249_add_4_5 .INJECT1_0 = "NO";
    defparam \genblk1.clock_cnt_2249_add_4_5 .INJECT1_1 = "NO";
    PFUMX mux_70_i5 (.BLUT(n4962[2]), .ALUT(n324[4]), .C0(n36490), .Z(SPI_DAT_O_31__N_4307[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;
    PFUMX mux_70_i4 (.BLUT(n4962[1]), .ALUT(n324[3]), .C0(n36490), .Z(SPI_DAT_O_31__N_4307[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;
    LUT4 mux_70_i21_4_lut (.A(reg_txdata[20]), .B(reg_rxdata[20]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i21_4_lut.init = 16'hcac0;
    CCU2C \genblk1.clock_cnt_2249_add_4_3  (.A0(\genblk1.clock_cnt [1]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(\genblk1.clock_cnt [2]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n27510), .COUT(n27511), .S0(n69[1]), 
          .S1(n69[2]));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249_add_4_3 .INIT0 = 16'haaa0;
    defparam \genblk1.clock_cnt_2249_add_4_3 .INIT1 = 16'haaa0;
    defparam \genblk1.clock_cnt_2249_add_4_3 .INJECT1_0 = "NO";
    defparam \genblk1.clock_cnt_2249_add_4_3 .INJECT1_1 = "NO";
    CCU2C \genblk1.clock_cnt_2249_add_4_1  (.A0(GND_net), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(\genblk1.clock_cnt [0]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .COUT(n27510), .S1(n69[0]));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249_add_4_1 .INIT0 = 16'h0000;
    defparam \genblk1.clock_cnt_2249_add_4_1 .INIT1 = 16'h555f;
    defparam \genblk1.clock_cnt_2249_add_4_1 .INJECT1_0 = "NO";
    defparam \genblk1.clock_cnt_2249_add_4_1 .INJECT1_1 = "NO";
    FD1S3DX latch_s_data_i1 (.D(n41329), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i1.GSR = "ENABLED";
    FD1S3DX latch_s_data_i2 (.D(n41330), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i2.GSR = "ENABLED";
    FD1S3DX latch_s_data_i3 (.D(n41331), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i3.GSR = "ENABLED";
    FD1S3DX latch_s_data_i4 (.D(n41332), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i4.GSR = "ENABLED";
    FD1S3DX latch_s_data_i5 (.D(n41333), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i5.GSR = "ENABLED";
    FD1S3DX latch_s_data_i6 (.D(n41334), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i6.GSR = "ENABLED";
    FD1S3DX latch_s_data_i7 (.D(n41335), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i7.GSR = "ENABLED";
    FD1S3DX latch_s_data_i8 (.D(\SHAREDBUS_DAT_I[8] ), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i8.GSR = "ENABLED";
    FD1S3DX latch_s_data_i9 (.D(\SHAREDBUS_DAT_I[9] ), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i9.GSR = "ENABLED";
    FD1S3DX latch_s_data_i10 (.D(\SHAREDBUS_DAT_I[10] ), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(latch_s_data[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i10.GSR = "ENABLED";
    FD1S3DX latch_s_data_i11 (.D(\SHAREDBUS_DAT_I[11] ), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(latch_s_data[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i11.GSR = "ENABLED";
    FD1S3DX latch_s_data_i12 (.D(\SHAREDBUS_DAT_I[12] ), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(latch_s_data[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i12.GSR = "ENABLED";
    FD1S3DX latch_s_data_i13 (.D(\SHAREDBUS_DAT_I[13] ), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(latch_s_data[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i13.GSR = "ENABLED";
    FD1S3DX latch_s_data_i14 (.D(\SHAREDBUS_DAT_I[14] ), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(latch_s_data[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i14.GSR = "ENABLED";
    FD1S3DX latch_s_data_i15 (.D(\SHAREDBUS_DAT_I[15] ), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(latch_s_data[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i15.GSR = "ENABLED";
    FD1S3DX latch_s_data_i16 (.D(n41336), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i16.GSR = "ENABLED";
    FD1S3DX latch_s_data_i17 (.D(n41337), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i17.GSR = "ENABLED";
    FD1S3DX latch_s_data_i18 (.D(n41338), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i18.GSR = "ENABLED";
    FD1S3DX latch_s_data_i19 (.D(n41339), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i19.GSR = "ENABLED";
    FD1S3DX latch_s_data_i20 (.D(n41340), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i20.GSR = "ENABLED";
    FD1S3DX latch_s_data_i21 (.D(n41341), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i21.GSR = "ENABLED";
    FD1S3DX latch_s_data_i22 (.D(n41342), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i22.GSR = "ENABLED";
    FD1S3DX latch_s_data_i23 (.D(n41343), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(latch_s_data[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i23.GSR = "ENABLED";
    FD1S3DX latch_s_data_i24 (.D(\SHAREDBUS_DAT_I[24] ), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(latch_s_data[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i24.GSR = "ENABLED";
    FD1S3DX latch_s_data_i25 (.D(\SHAREDBUS_DAT_I[25] ), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(latch_s_data[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i25.GSR = "ENABLED";
    FD1S3DX latch_s_data_i26 (.D(\SHAREDBUS_DAT_I[26] ), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(latch_s_data[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i26.GSR = "ENABLED";
    FD1S3DX latch_s_data_i27 (.D(\SHAREDBUS_DAT_I[27] ), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(latch_s_data[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i27.GSR = "ENABLED";
    FD1S3DX latch_s_data_i28 (.D(\SHAREDBUS_DAT_I[28] ), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(latch_s_data[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i28.GSR = "ENABLED";
    FD1S3DX latch_s_data_i29 (.D(\SHAREDBUS_DAT_I[29] ), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(latch_s_data[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i29.GSR = "ENABLED";
    FD1S3DX latch_s_data_i30 (.D(\SHAREDBUS_DAT_I[30] ), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(latch_s_data[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i30.GSR = "ENABLED";
    FD1S3DX latch_s_data_i31 (.D(\SHAREDBUS_DAT_I[31] ), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(latch_s_data[31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(201[8:41])
    defparam latch_s_data_i31.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i1 (.D(rx_shift_data[0]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i1.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i2 (.D(rx_shift_data[1]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i2.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i3 (.D(rx_shift_data[2]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i3.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i4 (.D(rx_shift_data[3]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i4.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i5 (.D(rx_shift_data[4]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i5.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i6 (.D(rx_shift_data[5]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i6.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i7 (.D(rx_shift_data[6]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i7.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i8 (.D(rx_shift_data[7]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i8.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i9 (.D(rx_shift_data[8]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i9.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i10 (.D(rx_shift_data[9]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i10.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i11 (.D(rx_shift_data[10]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i11.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i12 (.D(rx_shift_data[11]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i12.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i13 (.D(rx_shift_data[12]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i13.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i14 (.D(rx_shift_data[13]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i14.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i15 (.D(rx_shift_data[14]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i15.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i16 (.D(rx_shift_data[15]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i16.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i17 (.D(rx_shift_data[16]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i17.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i18 (.D(rx_shift_data[17]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i18.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i19 (.D(rx_shift_data[18]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i19.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i20 (.D(rx_shift_data[19]), .SP(REF_CLK_c_enable_1453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i20.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i21 (.D(rx_shift_data[20]), .SP(rx_shift_data_31__N_4339), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i21.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i22 (.D(rx_shift_data[21]), .SP(rx_shift_data_31__N_4339), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i22.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i23 (.D(rx_shift_data[22]), .SP(rx_shift_data_31__N_4339), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i23.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i24 (.D(rx_shift_data[23]), .SP(rx_shift_data_31__N_4339), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i24.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i25 (.D(rx_shift_data[24]), .SP(rx_shift_data_31__N_4339), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i25.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i26 (.D(rx_shift_data[25]), .SP(rx_shift_data_31__N_4339), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i26.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i27 (.D(rx_shift_data[26]), .SP(rx_shift_data_31__N_4339), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i27.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i28 (.D(rx_shift_data[27]), .SP(rx_shift_data_31__N_4339), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i28.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i29 (.D(rx_shift_data[28]), .SP(rx_shift_data_31__N_4339), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i29.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i30 (.D(rx_shift_data[29]), .SP(rx_shift_data_31__N_4339), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i30.GSR = "ENABLED";
    FD1P3DX rx_shift_data_i0_i31 (.D(rx_shift_data[30]), .SP(rx_shift_data_31__N_4339), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(rx_shift_data[31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(320[11] 325[9])
    defparam rx_shift_data_i0_i31.GSR = "ENABLED";
    FD1S3DX \genblk1.c_status_i1  (.D(\genblk1.n_status [1]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.c_status [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(349[10:31])
    defparam \genblk1.c_status_i1 .GSR = "ENABLED";
    FD1S3DX \genblk1.c_status_i2  (.D(\genblk1.n_status [2]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.c_status [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(349[10:31])
    defparam \genblk1.c_status_i2 .GSR = "ENABLED";
    FD1P3DX tx_shift_data_i1 (.D(tx_shift_data_31__N_4212[1]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i1.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i2 (.D(tx_shift_data_31__N_4212[2]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i2.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i3 (.D(tx_shift_data_31__N_4212[3]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i3.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i4 (.D(tx_shift_data_31__N_4212[4]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i4.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i5 (.D(tx_shift_data_31__N_4212[5]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i5.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i6 (.D(tx_shift_data_31__N_4212[6]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i6.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i7 (.D(tx_shift_data_31__N_4212[7]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i7.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i8 (.D(tx_shift_data_31__N_4212[8]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i8.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i9 (.D(tx_shift_data_31__N_4212[9]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i9.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i10 (.D(tx_shift_data_31__N_4212[10]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i10.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i11 (.D(tx_shift_data_31__N_4212[11]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i11.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i12 (.D(tx_shift_data_31__N_4212[12]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i12.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i13 (.D(tx_shift_data_31__N_4212[13]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i13.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i14 (.D(tx_shift_data_31__N_4212[14]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i14.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i15 (.D(tx_shift_data_31__N_4212[15]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i15.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i16 (.D(tx_shift_data_31__N_4212[16]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i16.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i17 (.D(tx_shift_data_31__N_4212[17]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i17.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i18 (.D(tx_shift_data_31__N_4212[18]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i18.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i19 (.D(tx_shift_data_31__N_4212[19]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i19.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i20 (.D(tx_shift_data_31__N_4212[20]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i20.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i21 (.D(tx_shift_data_31__N_4212[21]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i21.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i22 (.D(tx_shift_data_31__N_4212[22]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i22.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i23 (.D(tx_shift_data_31__N_4212[23]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i23.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i24 (.D(tx_shift_data_31__N_4212[24]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i24.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i25 (.D(tx_shift_data_31__N_4212[25]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i25.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i26 (.D(tx_shift_data_31__N_4212[26]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i26.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i27 (.D(tx_shift_data_31__N_4212[27]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i27.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i28 (.D(tx_shift_data_31__N_4212[28]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i28.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i29 (.D(tx_shift_data_31__N_4212[29]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i29.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i30 (.D(tx_shift_data_31__N_4212[30]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i30.GSR = "ENABLED";
    FD1P3DX tx_shift_data_i31 (.D(tx_shift_data_31__N_4212[31]), .SP(REF_CLK_c_enable_760), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(tx_shift_data[31])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam tx_shift_data_i31.GSR = "ENABLED";
    LUT4 mux_70_i20_4_lut (.A(reg_txdata[19]), .B(reg_rxdata[19]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i20_4_lut.init = 16'hcac0;
    LUT4 i25_4_lut (.A(\genblk1.c_status [2]), .B(\genblk1.c_status [1]), 
         .C(\genblk1.c_status [0]), .D(IO_SCK_c), .Z(n12)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B ((D)+!C)))) */ ;
    defparam i25_4_lut.init = 16'h6424;
    LUT4 i1_4_lut (.A(\genblk1.data_cnt [2]), .B(n35090), .C(\genblk1.data_cnt [3]), 
         .D(n11367), .Z(n15969)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut.init = 16'h0004;
    LUT4 i1_3_lut (.A(n12_adj_6337), .B(\genblk1.data_cnt [5]), .C(\genblk1.data_cnt [4]), 
         .Z(n35090)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i1_3_lut.init = 16'h0202;
    LUT4 mux_70_i19_4_lut (.A(reg_txdata[18]), .B(reg_rxdata[18]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i19_4_lut.init = 16'hcac0;
    LUT4 mux_70_i18_4_lut (.A(reg_txdata[17]), .B(reg_rxdata[17]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i18_4_lut.init = 16'hcac0;
    FD1P3DX \genblk1.data_cnt__i5  (.D(n12424), .SP(REF_CLK_c_enable_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\genblk1.data_cnt [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(402[12] 411[35])
    defparam \genblk1.data_cnt__i5 .GSR = "ENABLED";
    FD1P3DX \genblk1.data_cnt__i4  (.D(n12422), .SP(REF_CLK_c_enable_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\genblk1.data_cnt [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(402[12] 411[35])
    defparam \genblk1.data_cnt__i4 .GSR = "ENABLED";
    FD1P3DX \genblk1.data_cnt__i3  (.D(n28997), .SP(REF_CLK_c_enable_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\genblk1.data_cnt [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(402[12] 411[35])
    defparam \genblk1.data_cnt__i3 .GSR = "ENABLED";
    FD1P3DX \genblk1.data_cnt__i2  (.D(n12418), .SP(REF_CLK_c_enable_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\genblk1.data_cnt [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(402[12] 411[35])
    defparam \genblk1.data_cnt__i2 .GSR = "ENABLED";
    FD1P3DX \genblk1.data_cnt__i1  (.D(n9), .SP(REF_CLK_c_enable_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\genblk1.data_cnt [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(402[12] 411[35])
    defparam \genblk1.data_cnt__i1 .GSR = "ENABLED";
    LUT4 i3955_4_lut (.A(n35244), .B(\genblk1.n_status_2__N_4362 [1]), .C(\genblk1.c_status [0]), 
         .D(n29807), .Z(n9215)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i3955_4_lut.init = 16'h3035;
    LUT4 i6_3_lut (.A(n1), .B(reg_rxdata[0]), .C(dw00_cs), .Z(SPI_DAT_O_31__N_4307[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(140[28:35])
    defparam i6_3_lut.init = 16'hcaca;
    LUT4 i5_4_lut (.A(n35472), .B(reg_txdata[0]), .C(dw04_cs), .D(dw08_cs), 
         .Z(n1)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(140[28:35])
    defparam i5_4_lut.init = 16'hc0ca;
    LUT4 i1_3_lut_adj_717 (.A(dw0c_cs), .B(dw10_cs), .C(\genblk1.reg_ssmask [0]), 
         .Z(n35472)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(180[15] 186[9])
    defparam i1_3_lut_adj_717.init = 16'h4040;
    LUT4 i33280_3_lut_4_lut_rep_1145 (.A(\genblk1.c_status [1]), .B(n41383), 
         .C(IO_SCK_c), .D(n11367), .Z(n45179)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(431[17:38])
    defparam i33280_3_lut_4_lut_rep_1145.init = 16'h0002;
    LUT4 i33280_3_lut_4_lut_rep_1146 (.A(\genblk1.c_status [1]), .B(n41383), 
         .C(IO_SCK_c), .D(n11367), .Z(REF_CLK_c_enable_1453)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(431[17:38])
    defparam i33280_3_lut_4_lut_rep_1146.init = 16'h0002;
    LUT4 i1_3_lut_4_lut_adj_718 (.A(\genblk1.data_cnt [1]), .B(\genblk1.data_cnt [0]), 
         .C(\genblk1.data_cnt [2]), .D(n6264), .Z(n12418)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(411[22:34])
    defparam i1_3_lut_4_lut_adj_718.init = 16'h0078;
    LUT4 i1_3_lut_4_lut_adj_719 (.A(\genblk1.data_cnt [1]), .B(\genblk1.data_cnt [0]), 
         .C(\genblk1.data_cnt [3]), .D(\genblk1.data_cnt [2]), .Z(n7707)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(411[22:34])
    defparam i1_3_lut_4_lut_adj_719.init = 16'h8000;
    LUT4 i1_4_lut_adj_720 (.A(n41225), .B(\LM32D_ADR_O[1] ), .C(n41380), 
         .D(\LM32D_ADR_O[0] ), .Z(n30156)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_720.init = 16'hfaea;
    LUT4 i1_4_lut_adj_721 (.A(n41246), .B(n30986), .C(n41310), .D(n41304), 
         .Z(reg_wr_N_4472)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_4_lut_adj_721.init = 16'h2000;
    LUT4 i1_4_lut_adj_722 (.A(n41304), .B(n30986), .C(n41246), .D(n41310), 
         .Z(reg_rd_N_4474)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_722.init = 16'h1000;
    LUT4 i7006_4_lut (.A(\genblk1.c_status [1]), .B(n41442), .C(\genblk1.n_status_2__N_4368 [0]), 
         .D(n41383), .Z(n12376)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(277[11] 280[49])
    defparam i7006_4_lut.init = 16'hfcec;
    LUT4 i1_3_lut_adj_723 (.A(\genblk1.n_status [1]), .B(\genblk1.n_status [0]), 
         .C(\genblk1.n_status [2]), .Z(rx_latch_flag_N_4482)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_adj_723.init = 16'hf7f7;
    LUT4 i33377_3_lut (.A(\genblk1.n_status [0]), .B(\genblk1.n_status_2__N_4302 [0]), 
         .C(\genblk1.n_status_2__N_4305 ), .Z(\genblk1.n_status [0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(355[4] 397[11])
    defparam i33377_3_lut.init = 16'hcaca;
    LUT4 \genblk1.c_status_2__I_0_301_Mux_0_i7_3_lut  (.A(n3_adj_6338), .B(n6), 
         .C(\genblk1.c_status [2]), .Z(\genblk1.n_status_2__N_4302 [0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(357[8] 396[15])
    defparam \genblk1.c_status_2__I_0_301_Mux_0_i7_3_lut .init = 16'hcaca;
    LUT4 i14997_4_lut (.A(n35350), .B(\genblk1.c_status [1]), .C(n29807), 
         .D(\genblk1.c_status [0]), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(357[8] 396[15])
    defparam i14997_4_lut.init = 16'h3233;
    LUT4 i1_2_lut (.A(\genblk1.data_cnt [1]), .B(\genblk1.data_cnt [0]), 
         .Z(n35350)) /* synthesis lut_function=((B)+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[42:66])
    defparam i1_2_lut.init = 16'hdddd;
    LUT4 i1_4_lut_adj_724 (.A(\genblk1.data_cnt [2]), .B(n11367), .C(n35246), 
         .D(\genblk1.data_cnt [4]), .Z(n29807)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[42:66])
    defparam i1_4_lut_adj_724.init = 16'hfffe;
    LUT4 i1_2_lut_adj_725 (.A(\genblk1.data_cnt [3]), .B(\genblk1.data_cnt [5]), 
         .Z(n35246)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[42:66])
    defparam i1_2_lut_adj_725.init = 16'heeee;
    LUT4 i7004_4_lut (.A(reg_status_6__N_4260), .B(n41297), .C(reg_status[6]), 
         .D(rx_latch_flag_N_4482), .Z(n12374)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (C+!(D))+!B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(449[12] 452[24])
    defparam i7004_4_lut.init = 16'h50dc;
    LUT4 i7012_3_lut (.A(reg_status_7__N_4253), .B(reg_status_7__N_4251), 
         .C(reg_status[7]), .Z(n12382)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(466[12] 475[31])
    defparam i7012_3_lut.init = 16'hdcdc;
    LUT4 i1_3_lut_adj_726 (.A(dw00_cs), .B(reg_rd), .C(spiSPI_ACK_O), 
         .Z(reg_status_7__N_4253)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(473[16:46])
    defparam i1_3_lut_adj_726.init = 16'h8080;
    LUT4 i33140_4_lut (.A(\genblk1.n_status [2]), .B(n11367), .C(\genblk1.n_status [0]), 
         .D(\genblk1.n_status [1]), .Z(reg_status_7__N_4251)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(466[16:43])
    defparam i33140_4_lut.init = 16'h0002;
    LUT4 i15595_3_lut (.A(reg_status[7]), .B(reg_status_7__N_4253), .C(reg_status_7__N_4251), 
         .Z(REF_CLK_c_enable_74)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam i15595_3_lut.init = 16'hacac;
    LUT4 i33119_3_lut (.A(\genblk1.reg_ssmask [0]), .B(reg_control[10]), 
         .C(n12_adj_6339), .Z(SS_N_4105)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i33119_3_lut.init = 16'h5757;
    LUT4 i19_3_lut (.A(\genblk1.c_status [0]), .B(\genblk1.c_status [1]), 
         .C(\genblk1.c_status [2]), .Z(n12_adj_6339)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;
    defparam i19_3_lut.init = 16'h1c1c;
    LUT4 i1_2_lut_rep_978 (.A(\genblk1.c_status [2]), .B(\genblk1.c_status [0]), 
         .Z(n41383)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(349[10:31])
    defparam i1_2_lut_rep_978.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_892_3_lut (.A(\genblk1.c_status [2]), .B(\genblk1.c_status [0]), 
         .C(\genblk1.c_status [1]), .Z(n41297)) /* synthesis lut_function=(A+!(B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(349[10:31])
    defparam i1_2_lut_rep_892_3_lut.init = 16'hbfbf;
    LUT4 i1_2_lut_rep_804_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(\genblk1.c_status [0]), 
         .C(n11367), .D(\genblk1.c_status [1]), .Z(n41209)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(349[10:31])
    defparam i1_2_lut_rep_804_3_lut_4_lut.init = 16'hfbff;
    LUT4 SS_N_4113_I_0_2_lut_3_lut_4_lut (.A(\genblk1.c_status [2]), .B(\genblk1.c_status [0]), 
         .C(rx_latch_flag_N_4482), .D(\genblk1.c_status [1]), .Z(rx_latch_flag_N_4481)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(349[10:31])
    defparam SS_N_4113_I_0_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 reg_status_4__I_0_292_2_lut (.A(reg_status[4]), .B(reg_status[3]), 
         .Z(reg_status[8])) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(218[30:47])
    defparam reg_status_4__I_0_292_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_727 (.A(n35042), .B(n30986), .C(n41304), .D(read_wait_done), 
         .Z(n31773)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_727.init = 16'h2220;
    LUT4 i7_3_lut (.A(reg_txdata[8]), .B(reg_rxdata[8]), .C(dw00_cs), 
         .Z(n3)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(140[28:35])
    defparam i7_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_2_lut (.A(\genblk1.data_cnt [0]), .B(\genblk1.data_cnt [1]), 
         .Z(n35244)) /* synthesis lut_function=((B)+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(404[12] 411[35])
    defparam i1_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(\genblk1.data_cnt [0]), .B(\genblk1.c_status [2]), 
         .C(\genblk1.c_status [0]), .D(\genblk1.c_status [1]), .Z(n31971)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(404[12] 411[35])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i14571_2_lut_2_lut (.A(\genblk1.c_status [0]), .B(\genblk1.n_status_2__N_4368 [0]), 
         .Z(n1_adj_6340)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i14571_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_3_lut_3_lut (.A(\genblk1.c_status [2]), .B(\genblk1.c_status [1]), 
         .C(\genblk1.c_status [0]), .Z(n35456)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(404[12] 411[35])
    defparam i1_3_lut_3_lut.init = 16'h1414;
    LUT4 i1_4_lut_4_lut_4_lut (.A(\genblk1.c_status [2]), .B(\genblk1.c_status [1]), 
         .C(\genblk1.data_cnt [0]), .D(\genblk1.c_status [0]), .Z(n31905)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(404[12] 411[35])
    defparam i1_4_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i1_3_lut_rep_786_4_lut (.A(IO_SCK_c), .B(n41209), .C(\inst_reg[15] ), 
         .D(n10865), .Z(n41191)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_3_lut_rep_786_4_lut.init = 16'h0010;
    FD1S3DX \genblk1.clock_cnt_2249__i1  (.D(n87[1]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.clock_cnt [1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249__i1 .GSR = "ENABLED";
    FD1S3DX \genblk1.clock_cnt_2249__i2  (.D(n87[2]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.clock_cnt [2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249__i2 .GSR = "ENABLED";
    FD1S3DX \genblk1.clock_cnt_2249__i3  (.D(n87[3]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.clock_cnt [3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249__i3 .GSR = "ENABLED";
    FD1S3DX \genblk1.clock_cnt_2249__i4  (.D(n87[4]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.clock_cnt [4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249__i4 .GSR = "ENABLED";
    FD1S3DX \genblk1.clock_cnt_2249__i5  (.D(n87[5]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.clock_cnt [5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249__i5 .GSR = "ENABLED";
    FD1S3DX \genblk1.clock_cnt_2249__i6  (.D(n87[6]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.clock_cnt [6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249__i6 .GSR = "ENABLED";
    FD1S3DX \genblk1.clock_cnt_2249__i7  (.D(n87[7]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.clock_cnt [7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249__i7 .GSR = "ENABLED";
    FD1S3DX \genblk1.clock_cnt_2249__i8  (.D(n87[8]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.clock_cnt [8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249__i8 .GSR = "ENABLED";
    FD1S3DX \genblk1.clock_cnt_2249__i9  (.D(n87[9]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.clock_cnt [9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249__i9 .GSR = "ENABLED";
    FD1S3DX \genblk1.clock_cnt_2249__i10  (.D(n87[10]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.clock_cnt [10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249__i10 .GSR = "ENABLED";
    FD1S3DX \genblk1.clock_cnt_2249__i11  (.D(n87[11]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.clock_cnt [11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249__i11 .GSR = "ENABLED";
    FD1S3DX \genblk1.clock_cnt_2249__i12  (.D(n87[12]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.clock_cnt [12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249__i12 .GSR = "ENABLED";
    FD1S3DX \genblk1.clock_cnt_2249__i13  (.D(n87[13]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.clock_cnt [13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249__i13 .GSR = "ENABLED";
    FD1S3DX \genblk1.clock_cnt_2249__i14  (.D(n87[14]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.clock_cnt [14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249__i14 .GSR = "ENABLED";
    FD1S3DX \genblk1.clock_cnt_2249__i15  (.D(n87[15]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.clock_cnt [15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam \genblk1.clock_cnt_2249__i15 .GSR = "ENABLED";
    LUT4 i33328_2_lut (.A(n11393), .B(n11367), .Z(\genblk1.n_status_2__N_4362 [1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(343[23:36])
    defparam i33328_2_lut.init = 16'h2222;
    LUT4 i1_4_lut_adj_728 (.A(\genblk1.data_cnt [5]), .B(n41406), .C(n35254), 
         .D(\genblk1.data_cnt [3]), .Z(n11393)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_728.init = 16'h4000;
    LUT4 i1_2_lut_adj_729 (.A(\genblk1.data_cnt [4]), .B(IO_SCK_c), .Z(n35254)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_729.init = 16'h8888;
    LUT4 i33129_2_lut_3_lut_4_lut (.A(n41345), .B(n41344), .C(n30156), 
         .D(n41347), .Z(dw0c_cs_N_4470)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i33129_2_lut_3_lut_4_lut.init = 16'h0008;
    PFUMX i33568 (.BLUT(n38970), .ALUT(n38969), .C0(\genblk1.c_status [2]), 
          .Z(\genblk1.n_status [1]));
    LUT4 i14554_4_lut (.A(read_wait_done), .B(spiSPI_ACK_O), .C(n34742), 
         .D(n30986), .Z(n6364)) /* synthesis lut_function=(!(A (B)+!A (B+((D)+!C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(256[10] 259[30])
    defparam i14554_4_lut.init = 16'h2232;
    LUT4 reg_control_7__I_0_2_lut (.A(reg_control[7]), .B(reg_status[7]), 
         .Z(SPI_INT_O_N_4422)) /* synthesis lut_function=(A (B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(240[24:46])
    defparam reg_control_7__I_0_2_lut.init = 16'h8888;
    LUT4 reg_control_8__I_0_4_lut (.A(reg_control[8]), .B(reg_control[3]), 
         .C(SPI_INT_O_N_4420), .D(reg_status[3]), .Z(SPI_INT_O_N_4417)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(238[24:76])
    defparam reg_control_8__I_0_4_lut.init = 16'ha8a0;
    LUT4 reg_control_6__I_0_2_lut (.A(reg_control[6]), .B(reg_status[6]), 
         .Z(SPI_INT_O_N_4421)) /* synthesis lut_function=(A (B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(239[24:46])
    defparam reg_control_6__I_0_2_lut.init = 16'h8888;
    LUT4 reg_control_4__I_0_2_lut (.A(reg_control[4]), .B(reg_status[4]), 
         .Z(SPI_INT_O_N_4420)) /* synthesis lut_function=(A (B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(238[56:74])
    defparam reg_control_4__I_0_2_lut.init = 16'h8888;
    LUT4 i1_3_lut_rep_1001 (.A(\genblk1.data_cnt [1]), .B(\genblk1.data_cnt [0]), 
         .C(\genblk1.data_cnt [2]), .Z(n41406)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_rep_1001.init = 16'h8080;
    LUT4 i30534_2_lut_4_lut (.A(\genblk1.data_cnt [1]), .B(\genblk1.data_cnt [0]), 
         .C(\genblk1.data_cnt [2]), .D(\genblk1.data_cnt [3]), .Z(n28997)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;
    defparam i30534_2_lut_4_lut.init = 16'h7f80;
    LUT4 i33381_3_lut (.A(\genblk1.n_status [2]), .B(\genblk1.n_status_2__N_4302 [2]), 
         .C(\genblk1.n_status_2__N_4305 ), .Z(\genblk1.n_status [2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(355[4] 397[11])
    defparam i33381_3_lut.init = 16'hcaca;
    LUT4 \genblk1.c_status_2__I_0_301_Mux_2_i7_4_lut  (.A(n35354), .B(n6), 
         .C(\genblk1.c_status [2]), .D(\genblk1.n_status_2__N_4362 [1]), 
         .Z(\genblk1.n_status_2__N_4302 [2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(357[8] 396[15])
    defparam \genblk1.c_status_2__I_0_301_Mux_2_i7_4_lut .init = 16'hcac0;
    LUT4 i1_2_lut_adj_730 (.A(\genblk1.c_status [1]), .B(\genblk1.c_status [0]), 
         .Z(n35354)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_730.init = 16'h8888;
    LUT4 i33127_2_lut_3_lut_4_lut (.A(n41345), .B(n41344), .C(n30156), 
         .D(n41347), .Z(dw08_cs_N_4469)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(183[27:52])
    defparam i33127_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 reg_wr_I_0_288_2_lut (.A(reg_wr), .B(dw0c_cs), .Z(reg_control_10__N_4245)) /* synthesis lut_function=(A (B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(230[13:30])
    defparam reg_wr_I_0_288_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n41345), .B(n41344), .C(n953[0]), .D(n954[0]), 
         .Z(n34304)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(182[27:52])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hdfff;
    LUT4 i1_4_lut_adj_731 (.A(\genblk1.wait_one_tick_done ), .B(n6019), 
         .C(n41209), .D(IO_SCK_c), .Z(REF_CLK_c_enable_760)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(414[8:26])
    defparam i1_4_lut_adj_731.init = 16'hcecc;
    LUT4 i3968_3_lut (.A(tx_shift_data[31]), .B(reg_txdata[31]), .C(n6019), 
         .Z(n9228)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(430[12] 443[16])
    defparam i3968_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_732 (.A(n35456), .B(\genblk1.n_status [2]), .C(\genblk1.n_status [1]), 
         .D(\genblk1.n_status [0]), .Z(n6019)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_4_lut_adj_732.init = 16'h2000;
    LUT4 i33194_2_lut (.A(dw00_cs), .B(dw04_cs), .Z(n36490)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam i33194_2_lut.init = 16'heeee;
    LUT4 reg_wr_I_0_285_2_lut (.A(reg_wr), .B(dw10_cs), .Z(\genblk1.reg_ssmask_0__N_4110 )) /* synthesis lut_function=(A (B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(296[15:32])
    defparam reg_wr_I_0_285_2_lut.init = 16'h8888;
    LUT4 i33124_2_lut_3_lut_4_lut (.A(n41345), .B(n41344), .C(n30156), 
         .D(n41347), .Z(dw04_cs_N_4468)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(182[27:52])
    defparam i33124_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 mux_70_i17_4_lut (.A(reg_txdata[16]), .B(reg_rxdata[16]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i17_4_lut.init = 16'hcac0;
    LUT4 mux_70_i16_4_lut (.A(reg_txdata[15]), .B(reg_rxdata[15]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i16_4_lut.init = 16'hcac0;
    LUT4 mux_70_i15_4_lut (.A(reg_txdata[14]), .B(reg_rxdata[14]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i15_4_lut.init = 16'hcac0;
    LUT4 mux_70_i14_4_lut (.A(reg_txdata[13]), .B(reg_rxdata[13]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i14_4_lut.init = 16'hcac0;
    LUT4 mux_70_i13_4_lut (.A(reg_txdata[12]), .B(reg_rxdata[12]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i13_4_lut.init = 16'hcac0;
    LUT4 mux_70_i12_4_lut (.A(reg_txdata[11]), .B(reg_rxdata[11]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i12_4_lut.init = 16'hcac0;
    LUT4 i10_3_lut (.A(n5), .B(reg_rxdata[10]), .C(dw00_cs), .Z(SPI_DAT_O_31__N_4307[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(140[28:35])
    defparam i10_3_lut.init = 16'hcaca;
    LUT4 i9_4_lut (.A(n35468), .B(reg_txdata[10]), .C(dw04_cs), .D(dw08_cs), 
         .Z(n5)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(140[28:35])
    defparam i9_4_lut.init = 16'hc0ca;
    LUT4 i1_2_lut_adj_733 (.A(dw0c_cs), .B(reg_control[10]), .Z(n35468)) /* synthesis lut_function=(A (B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(180[15] 186[9])
    defparam i1_2_lut_adj_733.init = 16'h8888;
    LUT4 mux_70_i10_4_lut (.A(reg_txdata[9]), .B(reg_rxdata[9]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i10_4_lut.init = 16'hcac0;
    LUT4 mux_70_i6_3_lut (.A(n324[5]), .B(reg_rxdata[5]), .C(dw00_cs), 
         .Z(SPI_DAT_O_31__N_4307[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i6_3_lut.init = 16'hcaca;
    LUT4 mux_69_i6_4_lut (.A(dw08_cs), .B(reg_txdata[5]), .C(dw04_cs), 
         .D(reg_status[5]), .Z(n324[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(287[32] 291[47])
    defparam mux_69_i6_4_lut.init = 16'hcac0;
    LUT4 mux_70_i3_4_lut (.A(reg_txdata[2]), .B(reg_rxdata[2]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i3_4_lut.init = 16'hcac0;
    LUT4 mux_70_i2_4_lut (.A(reg_txdata[1]), .B(reg_rxdata[1]), .C(dw00_cs), 
         .D(dw04_cs), .Z(SPI_DAT_O_31__N_4307[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(286[32] 291[47])
    defparam mux_70_i2_4_lut.init = 16'hcac0;
    LUT4 i32521_3_lut_4_lut (.A(reg_control[8]), .B(dw0c_cs), .C(dw08_cs), 
         .D(reg_status[8]), .Z(n17939)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(289[32] 291[47])
    defparam i32521_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_adj_734 (.A(n6019), .B(reg_txdata[0]), .Z(tx_shift_data_31__N_4212[1])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_734.init = 16'h8888;
    LUT4 tx_shift_data_31__I_0_i3_3_lut (.A(tx_shift_data[1]), .B(reg_txdata[1]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i4_3_lut (.A(tx_shift_data[2]), .B(reg_txdata[2]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i5_3_lut (.A(tx_shift_data[3]), .B(reg_txdata[3]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i6_3_lut (.A(tx_shift_data[4]), .B(reg_txdata[4]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i7_3_lut (.A(tx_shift_data[5]), .B(reg_txdata[5]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i8_3_lut (.A(tx_shift_data[6]), .B(reg_txdata[6]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i9_3_lut (.A(tx_shift_data[7]), .B(reg_txdata[7]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i10_3_lut (.A(tx_shift_data[8]), .B(reg_txdata[8]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i11_3_lut (.A(tx_shift_data[9]), .B(reg_txdata[9]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i12_3_lut (.A(tx_shift_data[10]), .B(reg_txdata[10]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i13_3_lut (.A(tx_shift_data[11]), .B(reg_txdata[11]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i13_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i14_3_lut (.A(tx_shift_data[12]), .B(reg_txdata[12]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i14_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i15_3_lut (.A(tx_shift_data[13]), .B(reg_txdata[13]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i15_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i16_3_lut (.A(tx_shift_data[14]), .B(reg_txdata[14]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i16_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i17_3_lut (.A(tx_shift_data[15]), .B(reg_txdata[15]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i17_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i18_3_lut (.A(tx_shift_data[16]), .B(reg_txdata[16]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i18_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i19_3_lut (.A(tx_shift_data[17]), .B(reg_txdata[17]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i19_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i20_3_lut (.A(tx_shift_data[18]), .B(reg_txdata[18]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i20_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i21_3_lut (.A(tx_shift_data[19]), .B(reg_txdata[19]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i21_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i22_3_lut (.A(tx_shift_data[20]), .B(reg_txdata[20]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i22_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i23_3_lut (.A(tx_shift_data[21]), .B(reg_txdata[21]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i23_3_lut.init = 16'hcaca;
    LUT4 mux_69_i4_3_lut (.A(reg_txdata[3]), .B(reg_rxdata[3]), .C(dw00_cs), 
         .Z(n324[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(287[32] 291[47])
    defparam mux_69_i4_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i24_3_lut (.A(tx_shift_data[22]), .B(reg_txdata[22]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i24_3_lut.init = 16'hcaca;
    LUT4 i12634_4_lut (.A(reg_control[3]), .B(reg_status[3]), .C(dw08_cs), 
         .D(dw0c_cs), .Z(n4962[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(141[28:35])
    defparam i12634_4_lut.init = 16'hcac0;
    LUT4 tx_shift_data_31__I_0_i25_3_lut (.A(tx_shift_data[23]), .B(reg_txdata[23]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i25_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i26_3_lut (.A(tx_shift_data[24]), .B(reg_txdata[24]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i26_3_lut.init = 16'hcaca;
    LUT4 mux_69_i5_3_lut (.A(reg_txdata[4]), .B(reg_rxdata[4]), .C(dw00_cs), 
         .Z(n324[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(287[32] 291[47])
    defparam mux_69_i5_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i27_3_lut (.A(tx_shift_data[25]), .B(reg_txdata[25]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1662_i3_4_lut (.A(reg_control[4]), .B(reg_status[4]), .C(dw08_cs), 
         .D(dw0c_cs), .Z(n4962[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(288[32] 291[47])
    defparam mux_1662_i3_4_lut.init = 16'hcac0;
    LUT4 tx_shift_data_31__I_0_i28_3_lut (.A(tx_shift_data[26]), .B(reg_txdata[26]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i28_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i29_3_lut (.A(tx_shift_data[27]), .B(reg_txdata[27]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i29_3_lut.init = 16'hcaca;
    LUT4 mux_69_i7_3_lut (.A(reg_txdata[6]), .B(reg_rxdata[6]), .C(dw00_cs), 
         .Z(n324[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(287[32] 291[47])
    defparam mux_69_i7_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i30_3_lut (.A(tx_shift_data[28]), .B(reg_txdata[28]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1662_i5_4_lut (.A(reg_control[6]), .B(reg_status[6]), .C(dw08_cs), 
         .D(dw0c_cs), .Z(n4962[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(288[32] 291[47])
    defparam mux_1662_i5_4_lut.init = 16'hcac0;
    LUT4 tx_shift_data_31__I_0_i31_3_lut (.A(tx_shift_data[29]), .B(reg_txdata[29]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i31_3_lut.init = 16'hcaca;
    LUT4 tx_shift_data_31__I_0_i32_3_lut (.A(tx_shift_data[30]), .B(reg_txdata[30]), 
         .C(n6019), .Z(tx_shift_data_31__N_4212[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(437[12] 443[16])
    defparam tx_shift_data_31__I_0_i32_3_lut.init = 16'hcaca;
    LUT4 mux_69_i8_3_lut (.A(reg_txdata[7]), .B(reg_rxdata[7]), .C(dw00_cs), 
         .Z(n324[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(287[32] 291[47])
    defparam mux_69_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1662_i6_4_lut (.A(reg_control[7]), .B(reg_status[7]), .C(dw08_cs), 
         .D(dw0c_cs), .Z(n4962[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(288[32] 291[47])
    defparam mux_1662_i6_4_lut.init = 16'hcac0;
    LUT4 i1_3_lut_4_lut_adj_735 (.A(spiSPI_ACK_O), .B(reg_wr), .C(n41422), 
         .D(dw08_cs), .Z(REF_CLK_c_enable_73)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(457[16:59])
    defparam i1_3_lut_4_lut_adj_735.init = 16'h8880;
    LUT4 i1_2_lut_rep_1017 (.A(reg_status[6]), .B(dw04_cs), .Z(n41422)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(457[16:59])
    defparam i1_2_lut_rep_1017.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_736 (.A(reg_status[6]), .B(dw04_cs), .C(reg_wr), 
         .D(spiSPI_ACK_O), .Z(reg_status_4__N_4268)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(457[16:59])
    defparam i1_2_lut_3_lut_4_lut_adj_736.init = 16'h4000;
    LUT4 i1_2_lut_rep_1018 (.A(\genblk1.c_status [0]), .B(\genblk1.c_status [1]), 
         .Z(n41423)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i1_2_lut_rep_1018.init = 16'heeee;
    LUT4 i2_3_lut_4_lut (.A(\genblk1.c_status [0]), .B(\genblk1.c_status [1]), 
         .C(\genblk1.c_status [2]), .D(n11367), .Z(\genblk1.n_status_2__N_4305 )) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i2_3_lut_4_lut.init = 16'hefff;
    LUT4 i33085_2_lut_3_lut_4_lut (.A(\genblk1.c_status [0]), .B(\genblk1.c_status [1]), 
         .C(\genblk1.n_status_2__N_4368 [0]), .D(\genblk1.c_status [2]), 
         .Z(reg_status_5__N_4266)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(304[66:93])
    defparam i33085_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 reg_wr_I_0_293_2_lut_rep_1037 (.A(reg_wr), .B(dw04_cs), .Z(n41442)) /* synthesis lut_function=(A (B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[15:32])
    defparam reg_wr_I_0_293_2_lut_rep_1037.init = 16'h8888;
    LUT4 reg_status_6__N_4261_I_0_2_lut_3_lut (.A(reg_wr), .B(dw04_cs), 
         .C(reg_status[6]), .Z(reg_txdata_31__N_4306)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[15:32])
    defparam reg_status_6__N_4261_I_0_2_lut_3_lut.init = 16'h8080;
    LUT4 reg_status_6__I_175_2_lut_3_lut (.A(reg_wr), .B(dw04_cs), .C(spiSPI_ACK_O), 
         .Z(reg_status_6__N_4260)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(214[15:32])
    defparam reg_status_6__I_175_2_lut_3_lut.init = 16'h8080;
    LUT4 i15_2_lut_3_lut_4_lut (.A(\genblk1.c_status [1]), .B(n41383), .C(IO_SCK_c), 
         .D(n11367), .Z(SCLK_MASTER_N_4428)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(431[17:38])
    defparam i15_2_lut_3_lut_4_lut.init = 16'hf0d2;
    LUT4 i1_4_lut_adj_737 (.A(n34628), .B(n34618), .C(n34620), .D(\genblk1.clock_cnt [0]), 
         .Z(n11367)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i1_4_lut_adj_737.init = 16'hfeff;
    LUT4 i1_4_lut_adj_738 (.A(\genblk1.clock_cnt [1]), .B(\genblk1.clock_cnt [8]), 
         .C(\genblk1.clock_cnt [3]), .D(\genblk1.clock_cnt [11]), .Z(n34628)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_738.init = 16'hfffd;
    LUT4 i1_4_lut_adj_739 (.A(\genblk1.clock_cnt [12]), .B(n34606), .C(n34610), 
         .D(\genblk1.clock_cnt [5]), .Z(n34618)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_739.init = 16'hfffe;
    LUT4 i1_4_lut_adj_740 (.A(\genblk1.clock_cnt [2]), .B(\genblk1.clock_cnt [15]), 
         .C(n34604), .D(\genblk1.clock_cnt [10]), .Z(n34620)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_740.init = 16'hfffd;
    LUT4 i1_2_lut_adj_741 (.A(\genblk1.clock_cnt [13]), .B(\genblk1.clock_cnt [4]), 
         .Z(n34606)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_741.init = 16'heeee;
    LUT4 i1_2_lut_adj_742 (.A(\genblk1.clock_cnt [14]), .B(\genblk1.clock_cnt [6]), 
         .Z(n34610)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_742.init = 16'heeee;
    LUT4 i1_2_lut_adj_743 (.A(\genblk1.clock_cnt [9]), .B(\genblk1.clock_cnt [7]), 
         .Z(n34604)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_743.init = 16'heeee;
    LUT4 i1_4_lut_adj_744 (.A(n6264), .B(\genblk1.data_cnt [5]), .C(\genblk1.data_cnt [4]), 
         .D(n7707), .Z(n12424)) /* synthesis lut_function=(!(A+(B (C (D))+!B !(C (D))))) */ ;
    defparam i1_4_lut_adj_744.init = 16'h1444;
    LUT4 i1_3_lut_adj_745 (.A(n6264), .B(\genblk1.data_cnt [4]), .C(n7707), 
         .Z(n12422)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;
    defparam i1_3_lut_adj_745.init = 16'h1414;
    LUT4 i33234_3_lut (.A(n15969), .B(\genblk1.data_cnt [0]), .C(\genblk1.data_cnt [1]), 
         .Z(n9)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;
    defparam i33234_3_lut.init = 16'h1414;
    PFUMX \genblk1.c_status_2__I_0_301_Mux_0_i3  (.BLUT(n1_adj_6340), .ALUT(n9215), 
          .C0(\genblk1.c_status [1]), .Z(n3_adj_6338)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;
    
endmodule
//
// Verilog Description of module \wb_ebr_ctrl(SIZE=32768) 
//

module \wb_ebr_ctrl(SIZE=32768)  (\genblk1.write_data_7__N_3573 , REF_CLK_c, 
            REF_CLK_c_enable_1606, n41324, VCC_net, ebrEBR_DAT_O, \genblk1.read_address[10] , 
            \genblk1.write_address[10] , n3700, n5386, n5085, n41345, 
            n3432, n41323, n41255, \genblk1.state[2] , GND_net, \genblk1.raw_hazard , 
            ebrEBR_ACK_O, \genblk1.write_data_23__N_3541 , \genblk1.write_data_23__N_3549 , 
            \genblk1.write_data_31__N_3525 , \genblk1.write_data_15__N_3557 , 
            n12390, LM32D_DAT_O, \genblk1.read_data[20] , \genblk1.EBR_SEL_I_d[2] , 
            \genblk1.EBR_DAT_I_d[9] , \genblk1.EBR_DAT_I_d[10] , \genblk1.EBR_DAT_I_d[11] , 
            \genblk1.EBR_DAT_I_d[12] , \genblk1.EBR_DAT_I_d[13] , \genblk1.EBR_DAT_I_d[14] , 
            \genblk1.EBR_DAT_I_d[15] , \genblk1.EBR_DAT_I_d[16] , \genblk1.EBR_DAT_I_d[17] , 
            \genblk1.EBR_DAT_I_d[18] , \genblk1.EBR_DAT_I_d[19] , \genblk1.EBR_DAT_I_d[21] , 
            \genblk1.EBR_DAT_I_d[22] , \genblk1.EBR_DAT_I_d[23] , \genblk1.EBR_DAT_I_d[25] , 
            \genblk1.EBR_DAT_I_d[26] , \genblk1.EBR_DAT_I_d[27] , \genblk1.EBR_DAT_I_d[28] , 
            \genblk1.EBR_DAT_I_d[29] , \genblk1.EBR_DAT_I_d[30] , \genblk1.EBR_DAT_I_d[31] , 
            \genblk1.EBR_SEL_I_d[1] , n41238, n41309, \genblk1.EBR_SEL_I_d[3] , 
            n41239, \genblk1.write_data_d[2] , \genblk1.write_data_d[3] , 
            \genblk1.write_data_d[4] , \genblk1.write_data_d[6] , \genblk1.write_data_d[7] , 
            \genblk1.write_data_d[9] , \genblk1.write_data_d[10] , \genblk1.write_data_d[11] , 
            \genblk1.write_data_d[12] , \genblk1.write_data_d[13] , \genblk1.write_data_d[14] , 
            \genblk1.write_data_d[15] , \genblk1.write_data_d[16] , \genblk1.write_data_d[17] , 
            \genblk1.write_data_d[18] , \genblk1.write_data_d[19] , \genblk1.write_data_d[20] , 
            \genblk1.write_data_d[21] , \genblk1.write_data_d[22] , \genblk1.write_data_d[23] , 
            \genblk1.write_data_d[24] , \genblk1.write_data_d[25] , \genblk1.write_data_d[26] , 
            \genblk1.write_data_d[27] , \genblk1.write_data_d[28] , \genblk1.write_data_d[29] , 
            \genblk1.write_data_d[30] , \genblk1.write_data_d[31] , n41461, 
            n10004, \genblk1.pmi_address[3] , n10006, \genblk1.pmi_address[4] , 
            n10008, \genblk1.pmi_address[5] , n41488, \genblk1.pmi_address[6] , 
            n10012, \genblk1.pmi_address[7] , n41485, \genblk1.pmi_address[8] , 
            n10016, \genblk1.pmi_address[9] , n10018, \genblk1.pmi_address[10] , 
            n41482, \genblk1.pmi_address[11] , n10022, \genblk1.pmi_address[12] , 
            n10024, \genblk1.pmi_address[13] , n10026, \genblk1.pmi_address[14] , 
            n10028, n41221, n19, n41304, n41321, n41195, n5, n35788, 
            n41298, n20000, n41300, n41299, \SHAREDBUS_ADR_I[10] , 
            n41310, n41301, \SHAREDBUS_ADR_I[7] , n41346, \SHAREDBUS_ADR_I[5] , 
            n41347, n41344, n6038, n15, n41259, n29, \SHAREDBUS_ADR_I[26] , 
            \genblk1.read_data[6] , n41268, n41273, n41242, n41237, 
            \genblk1.read_data[7] , n41246, \SHAREDBUS_ADR_I[31] , \SHAREDBUS_ADR_I[15] , 
            n41222, \genblk1.write_data_23__N_3549[7] , \genblk1.write_data_23__N_3549[6] , 
            \genblk1.write_data_23__N_3549[5] , \genblk1.write_data_23__N_3549[3] , 
            n35840, n41260, \SHAREDBUS_ADR_I[16] , \genblk1.write_data_23__N_3549[2] , 
            n11843, \LM32D_ADR_O[1] , n41380, n3485, n6034, n41292, 
            n19822, n11831, n41307, n41390, n41306, n33, n71, 
            n3486, \counter[2] , n76, n21, \genblk1.read_data[24] , 
            \genblk1.write_data_23__N_3549[1] , \genblk1.write_data_31__N_3533[7] , 
            \genblk1.write_data_31__N_3533[6] , \genblk1.write_data_31__N_3533[5] , 
            \genblk1.write_data_31__N_3533[4] , \genblk1.write_data_31__N_3533[3] , 
            \genblk1.read_data[2] , \genblk1.read_data[3] , \genblk1.write_data_31__N_3533[2] , 
            \genblk1.write_data_31__N_3533[1] , \genblk1.write_data_15__N_3565[7] , 
            \genblk1.write_data_15__N_3565[6] , \genblk1.write_data_15__N_3565[5] , 
            \genblk1.read_data[4] , \genblk1.write_data_15__N_3565[4] , 
            \genblk1.write_data_15__N_3565[3] , \genblk1.write_data_15__N_3565[2] , 
            \genblk1.write_data_15__N_3565[1] ) /* synthesis syn_module_defined=1 */ ;
    input [7:0]\genblk1.write_data_7__N_3573 ;
    input REF_CLK_c;
    output REF_CLK_c_enable_1606;
    input n41324;
    input VCC_net;
    output [31:0]ebrEBR_DAT_O;
    input \genblk1.read_address[10] ;
    input \genblk1.write_address[10] ;
    output n3700;
    output n5386;
    output n5085;
    input n41345;
    output n3432;
    input n41323;
    input n41255;
    output \genblk1.state[2] ;
    input GND_net;
    output \genblk1.raw_hazard ;
    output ebrEBR_ACK_O;
    input [7:0]\genblk1.write_data_23__N_3541 ;
    input [7:0]\genblk1.write_data_23__N_3549 ;
    input [7:0]\genblk1.write_data_31__N_3525 ;
    input [7:0]\genblk1.write_data_15__N_3557 ;
    input n12390;
    input [31:0]LM32D_DAT_O;
    input \genblk1.read_data[20] ;
    output \genblk1.EBR_SEL_I_d[2] ;
    output \genblk1.EBR_DAT_I_d[9] ;
    output \genblk1.EBR_DAT_I_d[10] ;
    output \genblk1.EBR_DAT_I_d[11] ;
    output \genblk1.EBR_DAT_I_d[12] ;
    output \genblk1.EBR_DAT_I_d[13] ;
    output \genblk1.EBR_DAT_I_d[14] ;
    output \genblk1.EBR_DAT_I_d[15] ;
    output \genblk1.EBR_DAT_I_d[16] ;
    output \genblk1.EBR_DAT_I_d[17] ;
    output \genblk1.EBR_DAT_I_d[18] ;
    output \genblk1.EBR_DAT_I_d[19] ;
    output \genblk1.EBR_DAT_I_d[21] ;
    output \genblk1.EBR_DAT_I_d[22] ;
    output \genblk1.EBR_DAT_I_d[23] ;
    output \genblk1.EBR_DAT_I_d[25] ;
    output \genblk1.EBR_DAT_I_d[26] ;
    output \genblk1.EBR_DAT_I_d[27] ;
    output \genblk1.EBR_DAT_I_d[28] ;
    output \genblk1.EBR_DAT_I_d[29] ;
    output \genblk1.EBR_DAT_I_d[30] ;
    output \genblk1.EBR_DAT_I_d[31] ;
    output \genblk1.EBR_SEL_I_d[1] ;
    input n41238;
    input n41309;
    output \genblk1.EBR_SEL_I_d[3] ;
    input n41239;
    output \genblk1.write_data_d[2] ;
    output \genblk1.write_data_d[3] ;
    output \genblk1.write_data_d[4] ;
    output \genblk1.write_data_d[6] ;
    output \genblk1.write_data_d[7] ;
    output \genblk1.write_data_d[9] ;
    output \genblk1.write_data_d[10] ;
    output \genblk1.write_data_d[11] ;
    output \genblk1.write_data_d[12] ;
    output \genblk1.write_data_d[13] ;
    output \genblk1.write_data_d[14] ;
    output \genblk1.write_data_d[15] ;
    output \genblk1.write_data_d[16] ;
    output \genblk1.write_data_d[17] ;
    output \genblk1.write_data_d[18] ;
    output \genblk1.write_data_d[19] ;
    output \genblk1.write_data_d[20] ;
    output \genblk1.write_data_d[21] ;
    output \genblk1.write_data_d[22] ;
    output \genblk1.write_data_d[23] ;
    output \genblk1.write_data_d[24] ;
    output \genblk1.write_data_d[25] ;
    output \genblk1.write_data_d[26] ;
    output \genblk1.write_data_d[27] ;
    output \genblk1.write_data_d[28] ;
    output \genblk1.write_data_d[29] ;
    output \genblk1.write_data_d[30] ;
    output \genblk1.write_data_d[31] ;
    input n41461;
    input n10004;
    output \genblk1.pmi_address[3] ;
    input n10006;
    output \genblk1.pmi_address[4] ;
    input n10008;
    output \genblk1.pmi_address[5] ;
    input n41488;
    output \genblk1.pmi_address[6] ;
    input n10012;
    output \genblk1.pmi_address[7] ;
    input n41485;
    output \genblk1.pmi_address[8] ;
    input n10016;
    output \genblk1.pmi_address[9] ;
    input n10018;
    output \genblk1.pmi_address[10] ;
    input n41482;
    output \genblk1.pmi_address[11] ;
    input n10022;
    output \genblk1.pmi_address[12] ;
    input n10024;
    output \genblk1.pmi_address[13] ;
    input n10026;
    output \genblk1.pmi_address[14] ;
    input n10028;
    input n41221;
    input n19;
    input n41304;
    output n41321;
    input n41195;
    input n5;
    input n35788;
    input n41298;
    output n20000;
    input n41300;
    input n41299;
    input \SHAREDBUS_ADR_I[10] ;
    input n41310;
    input n41301;
    input \SHAREDBUS_ADR_I[7] ;
    input n41346;
    input \SHAREDBUS_ADR_I[5] ;
    input n41347;
    input n41344;
    output n6038;
    input n15;
    input n41259;
    input n29;
    input \SHAREDBUS_ADR_I[26] ;
    input \genblk1.read_data[6] ;
    input n41268;
    input n41273;
    input n41242;
    input n41237;
    input \genblk1.read_data[7] ;
    input n41246;
    input \SHAREDBUS_ADR_I[31] ;
    input \SHAREDBUS_ADR_I[15] ;
    input n41222;
    input \genblk1.write_data_23__N_3549[7] ;
    input \genblk1.write_data_23__N_3549[6] ;
    input \genblk1.write_data_23__N_3549[5] ;
    input \genblk1.write_data_23__N_3549[3] ;
    input n35840;
    input n41260;
    input \SHAREDBUS_ADR_I[16] ;
    input \genblk1.write_data_23__N_3549[2] ;
    output n11843;
    input \LM32D_ADR_O[1] ;
    input n41380;
    output n3485;
    input n6034;
    input n41292;
    output n19822;
    input n11831;
    input n41307;
    input n41390;
    input n41306;
    input n33;
    input n71;
    output n3486;
    input \counter[2] ;
    input n76;
    input n21;
    input \genblk1.read_data[24] ;
    input \genblk1.write_data_23__N_3549[1] ;
    input \genblk1.write_data_31__N_3533[7] ;
    input \genblk1.write_data_31__N_3533[6] ;
    input \genblk1.write_data_31__N_3533[5] ;
    input \genblk1.write_data_31__N_3533[4] ;
    input \genblk1.write_data_31__N_3533[3] ;
    input \genblk1.read_data[2] ;
    input \genblk1.read_data[3] ;
    input \genblk1.write_data_31__N_3533[2] ;
    input \genblk1.write_data_31__N_3533[1] ;
    input \genblk1.write_data_15__N_3565[7] ;
    input \genblk1.write_data_15__N_3565[6] ;
    input \genblk1.write_data_15__N_3565[5] ;
    input \genblk1.read_data[4] ;
    input \genblk1.write_data_15__N_3565[4] ;
    input \genblk1.write_data_15__N_3565[3] ;
    input \genblk1.write_data_15__N_3565[2] ;
    input \genblk1.write_data_15__N_3565[1] ;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    wire [7:0]\genblk1.write_data_7__N_3581 ;
    
    wire n37897;
    wire [31:0]\genblk1.write_data ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(241[31:41])
    wire [3:0]\genblk1.EBR_SEL_I_d ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(249[16:27])
    
    wire \genblk1.write_enable ;
    wire [12:0]\genblk1.read_address ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(243[31:43])
    wire [12:0]\genblk1.write_address ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(243[45:58])
    
    wire \genblk1.read_enable ;
    wire [31:0]\genblk1.write_data_d ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(241[43:55])
    wire [14:0]\genblk1.pmi_address ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(242[31:42])
    
    wire n9452;
    wire [2:0]\genblk1.state ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(255[13:18])
    
    wire n41426, n29035, n27357, \genblk1.raw_hazard_nxt_N_3774 ;
    wire [31:0]\genblk1.read_data ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(245[31:40])
    
    wire \genblk1.EBR_ACK_O_nxt , \genblk1.raw_hazard_nxt , n37896, n27356;
    wire [7:0]\genblk1.write_data_31__N_3533 ;
    wire [7:0]\genblk1.write_data_15__N_3565 ;
    
    wire REF_CLK_c_enable_1224, n5308, n20740;
    wire [31:0]\genblk1.EBR_DAT_I_d ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(248[31:42])
    wire [7:0]\genblk1.write_data_23__N_3549_c ;
    
    wire n20057, n34806, n35870, n30121, n31897, n31757;
    wire [2:0]n8;
    
    wire n34786, n9, n6013, n37902, n35288, n9_adj_6336, n35268, 
        n35702, n27355, n31566, n37901, n37900, n37899, n37898;
    
    PFUMX \genblk1.write_data_7__I_0_i5  (.BLUT(\genblk1.write_data_7__N_3573 [4]), 
          .ALUT(\genblk1.write_data_7__N_3581 [4]), .C0(n37897), .Z(\genblk1.write_data [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;
    FD1S3IX \genblk1.EBR_SEL_I_d__i0  (.D(n41324), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.EBR_SEL_I_d [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_SEL_I_d__i0 .GSR = "ENABLED";
    pmi_ram_dpEhnonessen321381923213819211e08d7f pmi_ram_dpECP5Uhexnonespeedsyncenablenoreg3213819232138192 (.Data({\genblk1.write_data }), 
            .WrAddress({\genblk1.write_address [12:11], \genblk1.write_address[10] , 
            \genblk1.write_address [9:0]}), .RdAddress({\genblk1.read_address [12:11], 
            \genblk1.read_address[10] , \genblk1.read_address [9:0]}), .Q({ebrEBR_DAT_O}), 
            .WrClock(REF_CLK_c), .RdClock(REF_CLK_c), .WrClockEn(VCC_net), 
            .RdClockEn(\genblk1.read_enable ), .WE(\genblk1.write_enable ), 
            .Reset(REF_CLK_c_enable_1606)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(668[2] 682[36])
    defparam pmi_ram_dpECP5Uhexnonespeedsyncenablenoreg3213819232138192.module_type = "pmi_ram_dp";
    defparam pmi_ram_dpECP5Uhexnonespeedsyncenablenoreg3213819232138192.pmi_family = "ECP5U";
    defparam pmi_ram_dpECP5Uhexnonespeedsyncenablenoreg3213819232138192.pmi_init_file_format = "hex";
    defparam pmi_ram_dpECP5Uhexnonespeedsyncenablenoreg3213819232138192.pmi_init_file = "none";
    defparam pmi_ram_dpECP5Uhexnonespeedsyncenablenoreg3213819232138192.pmi_optimization = "speed";
    defparam pmi_ram_dpECP5Uhexnonespeedsyncenablenoreg3213819232138192.pmi_resetmode = "sync";
    defparam pmi_ram_dpECP5Uhexnonespeedsyncenablenoreg3213819232138192.pmi_gsr = "enable";
    defparam pmi_ram_dpECP5Uhexnonespeedsyncenablenoreg3213819232138192.pmi_regmode = "noreg";
    defparam pmi_ram_dpECP5Uhexnonespeedsyncenablenoreg3213819232138192.pmi_rd_data_width = 32;
    defparam pmi_ram_dpECP5Uhexnonespeedsyncenablenoreg3213819232138192.pmi_rd_addr_width = 13;
    defparam pmi_ram_dpECP5Uhexnonespeedsyncenablenoreg3213819232138192.pmi_rd_addr_depth = 8192;
    defparam pmi_ram_dpECP5Uhexnonespeedsyncenablenoreg3213819232138192.pmi_wr_data_width = 32;
    defparam pmi_ram_dpECP5Uhexnonespeedsyncenablenoreg3213819232138192.pmi_wr_addr_width = 13;
    defparam pmi_ram_dpECP5Uhexnonespeedsyncenablenoreg3213819232138192.pmi_wr_addr_depth = 8192;
    FD1S3IX \genblk1.write_data_d__i0  (.D(\genblk1.write_data [0]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i0 .GSR = "ENABLED";
    FD1S3IX \genblk1.pmi_address_i0  (.D(n9452), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.pmi_address [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.pmi_address_i0 .GSR = "ENABLED";
    PFUMX \genblk1.write_data_7__I_0_i4  (.BLUT(\genblk1.write_data_7__N_3573 [3]), 
          .ALUT(\genblk1.write_data_7__N_3581 [3]), .C0(n37897), .Z(\genblk1.write_data [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;
    PFUMX \genblk1.write_data_7__I_0_i3  (.BLUT(\genblk1.write_data_7__N_3573 [2]), 
          .ALUT(\genblk1.write_data_7__N_3581 [2]), .C0(n37897), .Z(\genblk1.write_data [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;
    LUT4 i14535_3_lut_4_lut (.A(\genblk1.state [1]), .B(n41426), .C(n3700), 
         .D(n5386), .Z(n5085)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B (C+(D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(309[14:32])
    defparam i14535_3_lut_4_lut.init = 16'h00e1;
    LUT4 i5296_3_lut_4_lut (.A(\genblk1.state [1]), .B(n41426), .C(\genblk1.pmi_address [2]), 
         .D(n41345), .Z(n3432)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(309[14:32])
    defparam i5296_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23_3_lut_4_lut (.A(n41323), .B(\genblk1.state [0]), .C(n41255), 
         .D(\genblk1.state[2] ), .Z(n29035)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A (B (D)+!B !((D)+!C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(259[5] 289[12])
    defparam i23_3_lut_4_lut.init = 16'hcc1a;
    CCU2C \genblk1.read_address_12__I_0_13  (.A0(\genblk1.write_address [1]), 
          .B0(\genblk1.read_address [1]), .C0(\genblk1.write_address [0]), 
          .D0(\genblk1.read_address [0]), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27357), .S1(\genblk1.raw_hazard_nxt_N_3774 ));
    defparam \genblk1.read_address_12__I_0_13 .INIT0 = 16'h9009;
    defparam \genblk1.read_address_12__I_0_13 .INIT1 = 16'h0000;
    defparam \genblk1.read_address_12__I_0_13 .INJECT1_0 = "YES";
    defparam \genblk1.read_address_12__I_0_13 .INJECT1_1 = "NO";
    LUT4 EBR_DAT_O_31__I_0_161_i9_3_lut (.A(ebrEBR_DAT_O[8]), .B(\genblk1.write_data_d [8]), 
         .C(\genblk1.raw_hazard ), .Z(\genblk1.read_data [8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(316[20:52])
    defparam EBR_DAT_O_31__I_0_161_i9_3_lut.init = 16'hcaca;
    PFUMX \genblk1.write_data_7__I_0_i2  (.BLUT(\genblk1.write_data_7__N_3573 [1]), 
          .ALUT(\genblk1.write_data_7__N_3581 [1]), .C0(n37897), .Z(\genblk1.write_data [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;
    FD1S3IX EBR_ACK_O_146 (.D(\genblk1.EBR_ACK_O_nxt ), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(ebrEBR_ACK_O)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam EBR_ACK_O_146.GSR = "ENABLED";
    FD1S3IX \genblk1.raw_hazard_152  (.D(\genblk1.raw_hazard_nxt ), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.raw_hazard )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.raw_hazard_152 .GSR = "ENABLED";
    PFUMX mux_1090_i1 (.BLUT(\genblk1.write_data_23__N_3541 [0]), .ALUT(\genblk1.write_data_23__N_3549 [0]), 
          .C0(n37896), .Z(\genblk1.write_data [16]));
    CCU2C \genblk1.read_address_12__I_0_12  (.A0(\genblk1.write_address [5]), 
          .B0(\genblk1.read_address [5]), .C0(\genblk1.write_address [4]), 
          .D0(\genblk1.read_address [4]), .A1(\genblk1.write_address [3]), 
          .B1(\genblk1.read_address [3]), .C1(\genblk1.write_address [2]), 
          .D1(\genblk1.read_address [2]), .CIN(n27356), .COUT(n27357));
    defparam \genblk1.read_address_12__I_0_12 .INIT0 = 16'h9009;
    defparam \genblk1.read_address_12__I_0_12 .INIT1 = 16'h9009;
    defparam \genblk1.read_address_12__I_0_12 .INJECT1_0 = "YES";
    defparam \genblk1.read_address_12__I_0_12 .INJECT1_1 = "YES";
    PFUMX mux_1092_i1 (.BLUT(\genblk1.write_data_31__N_3525 [0]), .ALUT(\genblk1.write_data_31__N_3533 [0]), 
          .C0(n37896), .Z(\genblk1.write_data [24]));
    PFUMX mux_1088_i1 (.BLUT(\genblk1.write_data_15__N_3557 [0]), .ALUT(\genblk1.write_data_15__N_3565 [0]), 
          .C0(n37896), .Z(\genblk1.write_data [8]));
    LUT4 EBR_DAT_O_31__I_0_161_i1_3_lut (.A(ebrEBR_DAT_O[0]), .B(\genblk1.write_data_d [0]), 
         .C(\genblk1.raw_hazard ), .Z(\genblk1.read_data [0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(316[20:52])
    defparam EBR_DAT_O_31__I_0_161_i1_3_lut.init = 16'hcaca;
    PFUMX \genblk1.write_data_7__I_0_i1  (.BLUT(\genblk1.write_data_7__N_3573 [0]), 
          .ALUT(\genblk1.write_data_7__N_3581 [0]), .C0(n37896), .Z(\genblk1.write_data [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;
    FD1P3IX \genblk1.state__i0  (.D(n20740), .SP(REF_CLK_c_enable_1224), 
            .CD(n5308), .CK(REF_CLK_c), .Q(\genblk1.state [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.state__i0 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i0  (.D(LM32D_DAT_O[0]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d [0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i0 .GSR = "ENABLED";
    LUT4 mux_1089_i5_3_lut (.A(\genblk1.read_data[20] ), .B(\genblk1.EBR_DAT_I_d [20]), 
         .C(\genblk1.EBR_SEL_I_d[2] ), .Z(\genblk1.write_data_23__N_3549_c [4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam mux_1089_i5_3_lut.init = 16'hcaca;
    FD1S3IX \genblk1.EBR_DAT_I_d__i1  (.D(LM32D_DAT_O[1]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i1 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i2  (.D(LM32D_DAT_O[2]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i2 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i3  (.D(LM32D_DAT_O[3]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d [3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i3 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i4  (.D(LM32D_DAT_O[4]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d [4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i4 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i5  (.D(LM32D_DAT_O[5]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i5 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i6  (.D(LM32D_DAT_O[6]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i6 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i7  (.D(LM32D_DAT_O[7]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i7 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i8  (.D(LM32D_DAT_O[8]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d [8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i8 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i9  (.D(LM32D_DAT_O[9]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[9] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i9 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i10  (.D(LM32D_DAT_O[10]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[10] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i10 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i11  (.D(LM32D_DAT_O[11]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[11] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i11 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i12  (.D(LM32D_DAT_O[12]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[12] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i12 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i13  (.D(LM32D_DAT_O[13]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[13] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i13 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i14  (.D(LM32D_DAT_O[14]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[14] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i14 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i15  (.D(LM32D_DAT_O[15]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[15] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i15 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i16  (.D(LM32D_DAT_O[16]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[16] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i16 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i17  (.D(LM32D_DAT_O[17]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[17] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i17 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i18  (.D(LM32D_DAT_O[18]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[18] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i18 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i19  (.D(LM32D_DAT_O[19]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[19] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i19 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i20  (.D(LM32D_DAT_O[20]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d [20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i20 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i21  (.D(LM32D_DAT_O[21]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[21] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i21 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i22  (.D(LM32D_DAT_O[22]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[22] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i22 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i23  (.D(LM32D_DAT_O[23]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[23] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i23 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i24  (.D(LM32D_DAT_O[24]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d [24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i24 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i25  (.D(LM32D_DAT_O[25]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[25] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i25 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i26  (.D(LM32D_DAT_O[26]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[26] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i26 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i27  (.D(LM32D_DAT_O[27]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[27] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i27 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i28  (.D(LM32D_DAT_O[28]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[28] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i28 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i29  (.D(LM32D_DAT_O[29]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[29] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i29 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i30  (.D(LM32D_DAT_O[30]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[30] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i30 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_DAT_I_d__i31  (.D(LM32D_DAT_O[31]), .CK(REF_CLK_c), 
            .CD(n12390), .Q(\genblk1.EBR_DAT_I_d[31] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_DAT_I_d__i31 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_SEL_I_d__i1  (.D(n41238), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.EBR_SEL_I_d[1] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_SEL_I_d__i1 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_SEL_I_d__i2  (.D(n41309), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.EBR_SEL_I_d[2] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_SEL_I_d__i2 .GSR = "ENABLED";
    FD1S3IX \genblk1.EBR_SEL_I_d__i3  (.D(n41239), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.EBR_SEL_I_d[3] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.EBR_SEL_I_d__i3 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i1  (.D(\genblk1.write_data [1]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i1 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i2  (.D(\genblk1.write_data [2]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[2] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i2 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i3  (.D(\genblk1.write_data [3]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[3] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i3 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i4  (.D(\genblk1.write_data [4]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[4] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i4 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i5  (.D(\genblk1.write_data [5]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i5 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i6  (.D(\genblk1.write_data [6]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[6] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i6 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i7  (.D(\genblk1.write_data [7]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[7] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i7 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i8  (.D(\genblk1.write_data [8]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d [8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i8 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i9  (.D(\genblk1.write_data [9]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[9] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i9 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i10  (.D(\genblk1.write_data [10]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[10] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i10 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i11  (.D(\genblk1.write_data [11]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[11] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i11 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i12  (.D(\genblk1.write_data [12]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[12] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i12 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i13  (.D(\genblk1.write_data [13]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[13] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i13 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i14  (.D(\genblk1.write_data [14]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[14] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i14 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i15  (.D(\genblk1.write_data [15]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[15] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i15 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i16  (.D(\genblk1.write_data [16]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[16] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i16 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i17  (.D(\genblk1.write_data [17]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[17] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i17 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i18  (.D(\genblk1.write_data [18]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[18] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i18 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i19  (.D(\genblk1.write_data [19]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[19] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i19 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i20  (.D(\genblk1.write_data [20]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[20] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i20 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i21  (.D(\genblk1.write_data [21]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[21] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i21 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i22  (.D(\genblk1.write_data [22]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[22] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i22 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i23  (.D(\genblk1.write_data [23]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[23] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i23 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i24  (.D(\genblk1.write_data [24]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[24] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i24 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i25  (.D(\genblk1.write_data [25]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[25] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i25 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i26  (.D(\genblk1.write_data [26]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[26] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i26 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i27  (.D(\genblk1.write_data [27]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[27] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i27 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i28  (.D(\genblk1.write_data [28]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[28] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i28 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i29  (.D(\genblk1.write_data [29]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[29] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i29 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i30  (.D(\genblk1.write_data [30]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[30] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i30 .GSR = "ENABLED";
    FD1S3IX \genblk1.write_data_d__i31  (.D(\genblk1.write_data [31]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.write_data_d[31] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.write_data_d__i31 .GSR = "ENABLED";
    FD1S3IX \genblk1.pmi_address_i1  (.D(n41461), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.pmi_address [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.pmi_address_i1 .GSR = "ENABLED";
    FD1S3IX \genblk1.pmi_address_i2  (.D(n10004), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.pmi_address [2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.pmi_address_i2 .GSR = "ENABLED";
    FD1S3IX \genblk1.pmi_address_i3  (.D(n10006), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.pmi_address[3] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.pmi_address_i3 .GSR = "ENABLED";
    FD1S3IX \genblk1.pmi_address_i4  (.D(n10008), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.pmi_address[4] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.pmi_address_i4 .GSR = "ENABLED";
    FD1S3IX \genblk1.pmi_address_i5  (.D(n41488), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.pmi_address[5] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.pmi_address_i5 .GSR = "ENABLED";
    FD1S3IX \genblk1.pmi_address_i6  (.D(n10012), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.pmi_address[6] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.pmi_address_i6 .GSR = "ENABLED";
    FD1S3IX \genblk1.pmi_address_i7  (.D(n41485), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.pmi_address[7] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.pmi_address_i7 .GSR = "ENABLED";
    FD1S3IX \genblk1.pmi_address_i8  (.D(n10016), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.pmi_address[8] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.pmi_address_i8 .GSR = "ENABLED";
    FD1S3IX \genblk1.pmi_address_i9  (.D(n10018), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.pmi_address[9] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.pmi_address_i9 .GSR = "ENABLED";
    FD1S3IX \genblk1.pmi_address_i10  (.D(n41482), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.pmi_address[10] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.pmi_address_i10 .GSR = "ENABLED";
    FD1S3IX \genblk1.pmi_address_i11  (.D(n10022), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.pmi_address[11] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.pmi_address_i11 .GSR = "ENABLED";
    FD1S3IX \genblk1.pmi_address_i12  (.D(n10024), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.pmi_address[12] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.pmi_address_i12 .GSR = "ENABLED";
    FD1S3IX \genblk1.pmi_address_i13  (.D(n10026), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.pmi_address[13] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.pmi_address_i13 .GSR = "ENABLED";
    FD1S3IX \genblk1.pmi_address_i14  (.D(n10028), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\genblk1.pmi_address[14] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.pmi_address_i14 .GSR = "ENABLED";
    LUT4 EBR_DAT_O_31__I_0_161_i6_3_lut (.A(ebrEBR_DAT_O[5]), .B(\genblk1.write_data_d [5]), 
         .C(\genblk1.raw_hazard ), .Z(\genblk1.read_data [5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(316[20:52])
    defparam EBR_DAT_O_31__I_0_161_i6_3_lut.init = 16'hcaca;
    LUT4 i15552_4_lut (.A(n5308), .B(n20057), .C(n41221), .D(\genblk1.state [0]), 
         .Z(REF_CLK_c_enable_1224)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C (D)))) */ ;
    defparam i15552_4_lut.init = 16'hfaee;
    LUT4 i14793_4_lut (.A(n34806), .B(\genblk1.state[2] ), .C(n35870), 
         .D(n19), .Z(n20057)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B)) */ ;
    defparam i14793_4_lut.init = 16'hccce;
    LUT4 i1_4_lut (.A(\genblk1.state[2] ), .B(n41304), .C(n30121), .D(n31897), 
         .Z(\genblk1.write_enable )) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(327[12] 336[50])
    defparam i1_4_lut.init = 16'hece0;
    LUT4 i2_4_lut (.A(n41321), .B(n41195), .C(n5), .D(n35788), .Z(n31897)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_4_lut.init = 16'h0010;
    LUT4 \genblk1.pmi_address_14__I_0_i13_3_lut  (.A(\genblk1.pmi_address[14] ), 
         .B(n41298), .C(n20000), .Z(\genblk1.read_address [12])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(372[3:52])
    defparam \genblk1.pmi_address_14__I_0_i13_3_lut .init = 16'hacac;
    LUT4 \genblk1.pmi_address_14__I_0_i12_3_lut  (.A(\genblk1.pmi_address[13] ), 
         .B(n41300), .C(n20000), .Z(\genblk1.read_address [11])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(372[3:52])
    defparam \genblk1.pmi_address_14__I_0_i12_3_lut .init = 16'hacac;
    LUT4 \genblk1.pmi_address_14__I_0_i10_3_lut  (.A(\genblk1.pmi_address[11] ), 
         .B(n41299), .C(n20000), .Z(\genblk1.read_address [9])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(372[3:52])
    defparam \genblk1.pmi_address_14__I_0_i10_3_lut .init = 16'hacac;
    LUT4 \genblk1.pmi_address_14__I_0_i9_3_lut  (.A(\genblk1.pmi_address[10] ), 
         .B(\SHAREDBUS_ADR_I[10] ), .C(n20000), .Z(\genblk1.read_address [8])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(372[3:52])
    defparam \genblk1.pmi_address_14__I_0_i9_3_lut .init = 16'hacac;
    LUT4 \genblk1.pmi_address_14__I_0_i8_3_lut  (.A(\genblk1.pmi_address[9] ), 
         .B(n41310), .C(n20000), .Z(\genblk1.read_address [7])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(372[3:52])
    defparam \genblk1.pmi_address_14__I_0_i8_3_lut .init = 16'hacac;
    LUT4 \genblk1.pmi_address_14__I_0_i7_3_lut  (.A(\genblk1.pmi_address[8] ), 
         .B(n41301), .C(n20000), .Z(\genblk1.read_address [6])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(372[3:52])
    defparam \genblk1.pmi_address_14__I_0_i7_3_lut .init = 16'hacac;
    LUT4 \genblk1.pmi_address_14__I_0_i6_3_lut  (.A(\genblk1.pmi_address[7] ), 
         .B(\SHAREDBUS_ADR_I[7] ), .C(n20000), .Z(\genblk1.read_address [5])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(372[3:52])
    defparam \genblk1.pmi_address_14__I_0_i6_3_lut .init = 16'hacac;
    LUT4 \genblk1.pmi_address_14__I_0_i5_3_lut  (.A(\genblk1.pmi_address[6] ), 
         .B(n41346), .C(n20000), .Z(\genblk1.read_address [4])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(372[3:52])
    defparam \genblk1.pmi_address_14__I_0_i5_3_lut .init = 16'hacac;
    LUT4 \genblk1.pmi_address_14__I_0_i4_3_lut  (.A(\genblk1.pmi_address[5] ), 
         .B(\SHAREDBUS_ADR_I[5] ), .C(n20000), .Z(\genblk1.read_address [3])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(372[3:52])
    defparam \genblk1.pmi_address_14__I_0_i4_3_lut .init = 16'hacac;
    LUT4 \genblk1.pmi_address_14__I_0_i3_3_lut  (.A(\genblk1.pmi_address[4] ), 
         .B(n41347), .C(n20000), .Z(\genblk1.read_address [2])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(372[3:52])
    defparam \genblk1.pmi_address_14__I_0_i3_3_lut .init = 16'hacac;
    LUT4 \genblk1.pmi_address_14__I_0_i2_3_lut  (.A(\genblk1.pmi_address[3] ), 
         .B(n41344), .C(n20000), .Z(\genblk1.read_address [1])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(372[3:52])
    defparam \genblk1.pmi_address_14__I_0_i2_3_lut .init = 16'hacac;
    LUT4 \genblk1.pmi_address_14__I_0_i1_3_lut  (.A(\genblk1.pmi_address [2]), 
         .B(n41345), .C(n20000), .Z(\genblk1.read_address [0])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(372[3:52])
    defparam \genblk1.pmi_address_14__I_0_i1_3_lut .init = 16'hacac;
    LUT4 mux_1093_i13_3_lut (.A(n41298), .B(\genblk1.pmi_address[14] ), 
         .C(n6038), .Z(\genblk1.write_address [12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam mux_1093_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1093_i12_3_lut (.A(n41300), .B(\genblk1.pmi_address[13] ), 
         .C(n6038), .Z(\genblk1.write_address [11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam mux_1093_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1093_i10_3_lut (.A(n41299), .B(\genblk1.pmi_address[11] ), 
         .C(n6038), .Z(\genblk1.write_address [9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam mux_1093_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1093_i9_3_lut (.A(\SHAREDBUS_ADR_I[10] ), .B(\genblk1.pmi_address[10] ), 
         .C(n6038), .Z(\genblk1.write_address [8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam mux_1093_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1093_i8_3_lut (.A(n41310), .B(\genblk1.pmi_address[9] ), .C(n6038), 
         .Z(\genblk1.write_address [7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam mux_1093_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1093_i7_3_lut (.A(n41301), .B(\genblk1.pmi_address[8] ), .C(n6038), 
         .Z(\genblk1.write_address [6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam mux_1093_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1093_i6_3_lut (.A(\SHAREDBUS_ADR_I[7] ), .B(\genblk1.pmi_address[7] ), 
         .C(n6038), .Z(\genblk1.write_address [5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam mux_1093_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1093_i5_3_lut (.A(n41346), .B(\genblk1.pmi_address[6] ), .C(n6038), 
         .Z(\genblk1.write_address [4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam mux_1093_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1093_i4_3_lut (.A(\SHAREDBUS_ADR_I[5] ), .B(\genblk1.pmi_address[5] ), 
         .C(n6038), .Z(\genblk1.write_address [3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam mux_1093_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1093_i3_3_lut (.A(n41347), .B(\genblk1.pmi_address[4] ), .C(n6038), 
         .Z(\genblk1.write_address [2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam mux_1093_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1093_i2_3_lut (.A(n41344), .B(\genblk1.pmi_address[3] ), .C(n6038), 
         .Z(\genblk1.write_address [1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam mux_1093_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1093_i1_3_lut (.A(n41345), .B(\genblk1.pmi_address [2]), .C(n6038), 
         .Z(\genblk1.write_address [0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam mux_1093_i1_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_706 (.A(n31757), .B(n41304), .C(n41321), .D(n15), 
         .Z(\genblk1.read_enable )) /* synthesis lut_function=(A+!(B (C+!(D)))) */ ;
    defparam i2_4_lut_adj_706.init = 16'hbfbb;
    LUT4 i2_4_lut_adj_707 (.A(\genblk1.raw_hazard_nxt_N_3774 ), .B(\genblk1.state [1]), 
         .C(\genblk1.state [0]), .D(\genblk1.state[2] ), .Z(n31757)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+!(D)))) */ ;
    defparam i2_4_lut_adj_707.init = 16'h1300;
    LUT4 i1_3_lut (.A(\genblk1.state[2] ), .B(\genblk1.state [0]), .C(\genblk1.state [1]), 
         .Z(n6038)) /* synthesis lut_function=(!((B (C)+!B !(C))+!A)) */ ;
    defparam i1_3_lut.init = 16'h2828;
    LUT4 i14736_3_lut (.A(\genblk1.state [1]), .B(\genblk1.state [0]), .C(\genblk1.state[2] ), 
         .Z(n20000)) /* synthesis lut_function=(A+!(B (C)+!B !(C))) */ ;
    defparam i14736_3_lut.init = 16'hbebe;
    FD1P3AX \genblk1.state__i2  (.D(n8[2]), .SP(REF_CLK_c_enable_1224), 
            .CK(REF_CLK_c), .Q(\genblk1.state[2] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.state__i2 .GSR = "ENABLED";
    FD1P3IX \genblk1.state__i1  (.D(n29035), .SP(REF_CLK_c_enable_1224), 
            .CD(n5308), .CK(REF_CLK_c), .Q(\genblk1.state [1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam \genblk1.state__i1 .GSR = "ENABLED";
    LUT4 i32338_2_lut (.A(\genblk1.state [0]), .B(\genblk1.state [1]), .Z(n30121)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(327[12] 336[50])
    defparam i32338_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_708 (.A(n41259), .B(n34786), .C(n29), .D(\SHAREDBUS_ADR_I[26] ), 
         .Z(n34806)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_708.init = 16'h0004;
    LUT4 \genblk1.read_data_7__I_0_i7_3_lut  (.A(\genblk1.read_data[6] ), 
         .B(\genblk1.EBR_DAT_I_d [6]), .C(\genblk1.EBR_SEL_I_d [0]), .Z(\genblk1.write_data_7__N_3581 [6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(347[10:62])
    defparam \genblk1.read_data_7__I_0_i7_3_lut .init = 16'hcaca;
    LUT4 i30708_4_lut (.A(n41268), .B(n41273), .C(n41242), .D(n41237), 
         .Z(n35870)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30708_4_lut.init = 16'hfffe;
    LUT4 \genblk1.read_data_7__I_0_i8_3_lut  (.A(\genblk1.read_data[7] ), 
         .B(\genblk1.EBR_DAT_I_d [7]), .C(\genblk1.EBR_SEL_I_d [0]), .Z(\genblk1.write_data_7__N_3581 [7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(347[10:62])
    defparam \genblk1.read_data_7__I_0_i8_3_lut .init = 16'hcaca;
    LUT4 i1_4_lut_adj_709 (.A(n41246), .B(\SHAREDBUS_ADR_I[31] ), .C(\SHAREDBUS_ADR_I[15] ), 
         .D(ebrEBR_ACK_O), .Z(n34786)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_4_lut_adj_709.init = 16'h0020;
    LUT4 mux_1367_i1_4_lut (.A(n9), .B(\genblk1.state [0]), .C(\genblk1.state[2] ), 
         .D(n41222), .Z(n20740)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(259[5] 289[12])
    defparam mux_1367_i1_4_lut.init = 16'h3530;
    PFUMX mux_1090_i8 (.BLUT(\genblk1.write_data_23__N_3541 [7]), .ALUT(\genblk1.write_data_23__N_3549[7] ), 
          .C0(n6013), .Z(\genblk1.write_data [23]));
    PFUMX mux_1090_i7 (.BLUT(\genblk1.write_data_23__N_3541 [6]), .ALUT(\genblk1.write_data_23__N_3549[6] ), 
          .C0(n6013), .Z(\genblk1.write_data [22]));
    PFUMX mux_1090_i6 (.BLUT(\genblk1.write_data_23__N_3541 [5]), .ALUT(\genblk1.write_data_23__N_3549[5] ), 
          .C0(n6013), .Z(\genblk1.write_data [21]));
    PFUMX mux_1090_i5 (.BLUT(\genblk1.write_data_23__N_3541 [4]), .ALUT(\genblk1.write_data_23__N_3549_c [4]), 
          .C0(n6013), .Z(\genblk1.write_data [20]));
    PFUMX mux_1090_i4 (.BLUT(\genblk1.write_data_23__N_3541 [3]), .ALUT(\genblk1.write_data_23__N_3549[3] ), 
          .C0(n37902), .Z(\genblk1.write_data [19]));
    LUT4 EBR_DAT_O_31__I_0_161_i2_3_lut (.A(ebrEBR_DAT_O[1]), .B(\genblk1.write_data_d [1]), 
         .C(\genblk1.raw_hazard ), .Z(\genblk1.read_data [1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(316[20:52])
    defparam EBR_DAT_O_31__I_0_161_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_710 (.A(n35288), .B(n9_adj_6336), .C(n35840), .D(n19), 
         .Z(\genblk1.EBR_ACK_O_nxt )) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_710.init = 16'hccce;
    LUT4 i1_4_lut_adj_711 (.A(n41260), .B(n35268), .C(n29), .D(\SHAREDBUS_ADR_I[16] ), 
         .Z(n35288)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_711.init = 16'h0004;
    LUT4 i1_4_lut_adj_712 (.A(n41246), .B(\SHAREDBUS_ADR_I[31] ), .C(\SHAREDBUS_ADR_I[15] ), 
         .D(n35702), .Z(n35268)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_4_lut_adj_712.init = 16'h0020;
    LUT4 i1_4_lut_adj_713 (.A(\genblk1.state [1]), .B(\genblk1.raw_hazard_nxt_N_3774 ), 
         .C(\genblk1.state[2] ), .D(\genblk1.state [0]), .Z(\genblk1.raw_hazard_nxt )) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_713.init = 16'h4000;
    PFUMX mux_1090_i3 (.BLUT(\genblk1.write_data_23__N_3541 [2]), .ALUT(\genblk1.write_data_23__N_3549[2] ), 
          .C0(n37902), .Z(\genblk1.write_data [18]));
    CCU2C \genblk1.read_address_12__I_0_10  (.A0(\genblk1.write_address [9]), 
          .B0(\genblk1.read_address [9]), .C0(\genblk1.write_address [8]), 
          .D0(\genblk1.read_address [8]), .A1(\genblk1.write_address [7]), 
          .B1(\genblk1.read_address [7]), .C1(\genblk1.write_address [6]), 
          .D1(\genblk1.read_address [6]), .CIN(n27355), .COUT(n27356));
    defparam \genblk1.read_address_12__I_0_10 .INIT0 = 16'h9009;
    defparam \genblk1.read_address_12__I_0_10 .INIT1 = 16'h9009;
    defparam \genblk1.read_address_12__I_0_10 .INJECT1_0 = "YES";
    defparam \genblk1.read_address_12__I_0_10 .INJECT1_1 = "YES";
    CCU2C \genblk1.read_address_12__I_0_0  (.A0(\genblk1.write_address [12]), 
          .B0(\genblk1.read_address [12]), .C0(GND_net), .D0(VCC_net), 
          .A1(\genblk1.write_address [11]), .B1(\genblk1.read_address [11]), 
          .C1(\genblk1.write_address[10] ), .D1(\genblk1.read_address[10] ), 
          .COUT(n27355));   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(295[30:61])
    defparam \genblk1.read_address_12__I_0_0 .INIT0 = 16'h0009;
    defparam \genblk1.read_address_12__I_0_0 .INIT1 = 16'h9009;
    defparam \genblk1.read_address_12__I_0_0 .INJECT1_0 = "NO";
    defparam \genblk1.read_address_12__I_0_0 .INJECT1_1 = "YES";
    LUT4 i1_2_lut (.A(\genblk1.state [0]), .B(\genblk1.state [1]), .Z(n11843)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(309[14:32])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i4643_4_lut (.A(\LM32D_ADR_O[1] ), .B(\genblk1.pmi_address [1]), 
         .C(n41321), .D(n41380), .Z(n3485)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(434[7] 442[10])
    defparam i4643_4_lut.init = 16'hcac0;
    LUT4 i1_4_lut_adj_714 (.A(n6034), .B(n41292), .C(n19822), .D(n41321), 
         .Z(n3700)) /* synthesis lut_function=(A (B (D))+!A !((C+(D))+!B)) */ ;
    defparam i1_4_lut_adj_714.init = 16'h8804;
    LUT4 i14558_4_lut (.A(n31566), .B(n11831), .C(n41309), .D(n41307), 
         .Z(n19822)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i14558_4_lut.init = 16'haaa8;
    LUT4 i1_4_lut_adj_715 (.A(n41390), .B(n41324), .C(n41306), .D(n33), 
         .Z(n31566)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(309[87:109])
    defparam i1_4_lut_adj_715.init = 16'hfefc;
    LUT4 mux_1222_i1_4_lut (.A(n41321), .B(\genblk1.pmi_address [0]), .C(n3700), 
         .D(n71), .Z(n3486)) /* synthesis lut_function=(A (B (C))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(434[7] 442[10])
    defparam mux_1222_i1_4_lut.init = 16'h8580;
    LUT4 i20_3_lut_4_lut (.A(n41304), .B(\counter[2] ), .C(n71), .D(n76), 
         .Z(n9452)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i20_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_3_lut_4_lut (.A(\counter[2] ), .B(n41304), .C(n6034), .D(n19822), 
         .Z(n5386)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h0200;
    LUT4 counter_2__I_0_1_lut_rep_1016 (.A(\counter[2] ), .Z(REF_CLK_c_enable_1606)) /* synthesis lut_function=(!(A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(466[18:29])
    defparam counter_2__I_0_1_lut_rep_1016.init = 16'h5555;
    LUT4 i1912_2_lut_2_lut (.A(\counter[2] ), .B(\genblk1.state [1]), .Z(n5308)) /* synthesis lut_function=((B)+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(466[18:29])
    defparam i1912_2_lut_2_lut.init = 16'hdddd;
    LUT4 i11_2_lut_4_lut (.A(n41390), .B(n33), .C(n21), .D(n41304), 
         .Z(n9)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(309[87:109])
    defparam i11_2_lut_4_lut.init = 16'h8a00;
    LUT4 i1_2_lut_rep_1021 (.A(\genblk1.state[2] ), .B(\genblk1.state [0]), 
         .Z(n41426)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(309[14:32])
    defparam i1_2_lut_rep_1021.init = 16'heeee;
    LUT4 i1_2_lut_3_lut (.A(\genblk1.state[2] ), .B(\genblk1.state [0]), 
         .C(\genblk1.state [1]), .Z(n9_adj_6336)) /* synthesis lut_function=(!(A (C)+!A ((C)+!B))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(309[14:32])
    defparam i1_2_lut_3_lut.init = 16'h0e0e;
    LUT4 i30543_2_lut_3_lut_4_lut (.A(\genblk1.state[2] ), .B(\genblk1.state [0]), 
         .C(ebrEBR_ACK_O), .D(\genblk1.state [1]), .Z(n35702)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(309[14:32])
    defparam i30543_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_916_3_lut (.A(\genblk1.state[2] ), .B(\genblk1.state [0]), 
         .C(\genblk1.state [1]), .Z(n41321)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(309[14:32])
    defparam i1_2_lut_rep_916_3_lut.init = 16'hfefe;
    LUT4 i1_rep_133_2_lut_3_lut (.A(\genblk1.state [1]), .B(\genblk1.state [0]), 
         .C(\genblk1.state[2] ), .Z(n37897)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_rep_133_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_rep_132_2_lut_3_lut (.A(\genblk1.state [1]), .B(\genblk1.state [0]), 
         .C(\genblk1.state[2] ), .Z(n37896)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_rep_132_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_3_lut_adj_716 (.A(\genblk1.state [1]), .B(\genblk1.state [0]), 
         .C(\genblk1.state[2] ), .Z(n6013)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut_adj_716.init = 16'h7070;
    LUT4 i1_rep_138_2_lut_3_lut (.A(\genblk1.state [1]), .B(\genblk1.state [0]), 
         .C(\genblk1.state[2] ), .Z(n37902)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_rep_138_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_rep_137_2_lut_3_lut (.A(\genblk1.state [1]), .B(\genblk1.state [0]), 
         .C(\genblk1.state[2] ), .Z(n37901)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_rep_137_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_rep_136_2_lut_3_lut (.A(\genblk1.state [1]), .B(\genblk1.state [0]), 
         .C(\genblk1.state[2] ), .Z(n37900)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_rep_136_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_rep_135_2_lut_3_lut (.A(\genblk1.state [1]), .B(\genblk1.state [0]), 
         .C(\genblk1.state[2] ), .Z(n37899)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_rep_135_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_rep_134_2_lut_3_lut (.A(\genblk1.state [1]), .B(\genblk1.state [0]), 
         .C(\genblk1.state[2] ), .Z(n37898)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_rep_134_2_lut_3_lut.init = 16'h7070;
    LUT4 \genblk1.read_data_7__I_0_i1_3_lut  (.A(\genblk1.read_data [0]), 
         .B(\genblk1.EBR_DAT_I_d [0]), .C(\genblk1.EBR_SEL_I_d [0]), .Z(\genblk1.write_data_7__N_3581 [0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(347[10:62])
    defparam \genblk1.read_data_7__I_0_i1_3_lut .init = 16'hcaca;
    LUT4 mux_1087_i1_3_lut (.A(\genblk1.read_data [8]), .B(\genblk1.EBR_DAT_I_d [8]), 
         .C(\genblk1.EBR_SEL_I_d[1] ), .Z(\genblk1.write_data_15__N_3565 [0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam mux_1087_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1091_i1_3_lut (.A(\genblk1.read_data[24] ), .B(\genblk1.EBR_DAT_I_d [24]), 
         .C(\genblk1.EBR_SEL_I_d[3] ), .Z(\genblk1.write_data_31__N_3533 [0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam mux_1091_i1_3_lut.init = 16'hcaca;
    PFUMX mux_1090_i2 (.BLUT(\genblk1.write_data_23__N_3541 [1]), .ALUT(\genblk1.write_data_23__N_3549[1] ), 
          .C0(n37902), .Z(\genblk1.write_data [17]));
    PFUMX mux_1092_i8 (.BLUT(\genblk1.write_data_31__N_3525 [7]), .ALUT(\genblk1.write_data_31__N_3533[7] ), 
          .C0(n37902), .Z(\genblk1.write_data [31]));
    PFUMX mux_1092_i7 (.BLUT(\genblk1.write_data_31__N_3525 [6]), .ALUT(\genblk1.write_data_31__N_3533[6] ), 
          .C0(n37901), .Z(\genblk1.write_data [30]));
    PFUMX mux_1092_i6 (.BLUT(\genblk1.write_data_31__N_3525 [5]), .ALUT(\genblk1.write_data_31__N_3533[5] ), 
          .C0(n37901), .Z(\genblk1.write_data [29]));
    LUT4 \genblk1.read_data_7__I_0_i2_3_lut  (.A(\genblk1.read_data [1]), 
         .B(\genblk1.EBR_DAT_I_d [1]), .C(\genblk1.EBR_SEL_I_d [0]), .Z(\genblk1.write_data_7__N_3581 [1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(347[10:62])
    defparam \genblk1.read_data_7__I_0_i2_3_lut .init = 16'hcaca;
    PFUMX mux_1092_i5 (.BLUT(\genblk1.write_data_31__N_3525 [4]), .ALUT(\genblk1.write_data_31__N_3533[4] ), 
          .C0(n37901), .Z(\genblk1.write_data [28]));
    PFUMX mux_1092_i4 (.BLUT(\genblk1.write_data_31__N_3525 [3]), .ALUT(\genblk1.write_data_31__N_3533[3] ), 
          .C0(n37901), .Z(\genblk1.write_data [27]));
    LUT4 \genblk1.read_data_7__I_0_i3_3_lut  (.A(\genblk1.read_data[2] ), 
         .B(\genblk1.EBR_DAT_I_d [2]), .C(\genblk1.EBR_SEL_I_d [0]), .Z(\genblk1.write_data_7__N_3581 [2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(347[10:62])
    defparam \genblk1.read_data_7__I_0_i3_3_lut .init = 16'hcaca;
    LUT4 \genblk1.read_data_7__I_0_i4_3_lut  (.A(\genblk1.read_data[3] ), 
         .B(\genblk1.EBR_DAT_I_d [3]), .C(\genblk1.EBR_SEL_I_d [0]), .Z(\genblk1.write_data_7__N_3581 [3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(347[10:62])
    defparam \genblk1.read_data_7__I_0_i4_3_lut .init = 16'hcaca;
    PFUMX mux_1092_i3 (.BLUT(\genblk1.write_data_31__N_3525 [2]), .ALUT(\genblk1.write_data_31__N_3533[2] ), 
          .C0(n37900), .Z(\genblk1.write_data [26]));
    PFUMX mux_1092_i2 (.BLUT(\genblk1.write_data_31__N_3525 [1]), .ALUT(\genblk1.write_data_31__N_3533[1] ), 
          .C0(n37900), .Z(\genblk1.write_data [25]));
    PFUMX mux_1088_i8 (.BLUT(\genblk1.write_data_15__N_3557 [7]), .ALUT(\genblk1.write_data_15__N_3565[7] ), 
          .C0(n37900), .Z(\genblk1.write_data [15]));
    PFUMX mux_1088_i7 (.BLUT(\genblk1.write_data_15__N_3557 [6]), .ALUT(\genblk1.write_data_15__N_3565[6] ), 
          .C0(n37900), .Z(\genblk1.write_data [14]));
    PFUMX mux_1088_i6 (.BLUT(\genblk1.write_data_15__N_3557 [5]), .ALUT(\genblk1.write_data_15__N_3565[5] ), 
          .C0(n37899), .Z(\genblk1.write_data [13]));
    LUT4 \genblk1.read_data_7__I_0_i5_3_lut  (.A(\genblk1.read_data[4] ), 
         .B(\genblk1.EBR_DAT_I_d [4]), .C(\genblk1.EBR_SEL_I_d [0]), .Z(\genblk1.write_data_7__N_3581 [4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(347[10:62])
    defparam \genblk1.read_data_7__I_0_i5_3_lut .init = 16'hcaca;
    PFUMX mux_1088_i5 (.BLUT(\genblk1.write_data_15__N_3557 [4]), .ALUT(\genblk1.write_data_15__N_3565[4] ), 
          .C0(n37899), .Z(\genblk1.write_data [12]));
    LUT4 \genblk1.read_data_7__I_0_i6_3_lut  (.A(\genblk1.read_data [5]), 
         .B(\genblk1.EBR_DAT_I_d [5]), .C(\genblk1.EBR_SEL_I_d [0]), .Z(\genblk1.write_data_7__N_3581 [5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(347[10:62])
    defparam \genblk1.read_data_7__I_0_i6_3_lut .init = 16'hcaca;
    PFUMX mux_1088_i4 (.BLUT(\genblk1.write_data_15__N_3557 [3]), .ALUT(\genblk1.write_data_15__N_3565[3] ), 
          .C0(n37899), .Z(\genblk1.write_data [11]));
    PFUMX mux_1088_i3 (.BLUT(\genblk1.write_data_15__N_3557 [2]), .ALUT(\genblk1.write_data_15__N_3565[2] ), 
          .C0(n37899), .Z(\genblk1.write_data [10]));
    PFUMX mux_1088_i2 (.BLUT(\genblk1.write_data_15__N_3557 [1]), .ALUT(\genblk1.write_data_15__N_3565[1] ), 
          .C0(n37898), .Z(\genblk1.write_data [9]));
    PFUMX \genblk1.write_data_7__I_0_i8  (.BLUT(\genblk1.write_data_7__N_3573 [7]), 
          .ALUT(\genblk1.write_data_7__N_3581 [7]), .C0(n37898), .Z(\genblk1.write_data [7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;
    LUT4 i15150_4_lut (.A(n9), .B(n5308), .C(\genblk1.state[2] ), .D(n41222), 
         .Z(n8[2])) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/wb_ebr_ctrl/rtl/verilog/wb_ebr_ctrl.v(422[10] 442[10])
    defparam i15150_4_lut.init = 16'h3230;
    PFUMX \genblk1.write_data_7__I_0_i7  (.BLUT(\genblk1.write_data_7__N_3573 [6]), 
          .ALUT(\genblk1.write_data_7__N_3581 [6]), .C0(n37898), .Z(\genblk1.write_data [6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;
    PFUMX \genblk1.write_data_7__I_0_i6  (.BLUT(\genblk1.write_data_7__N_3573 [5]), 
          .ALUT(\genblk1.write_data_7__N_3581 [5]), .C0(n37898), .Z(\genblk1.write_data [5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=668, LSE_RLINE=682 */ ;
    
endmodule
//
// Verilog Description of module arbiter2
//

module arbiter2 (LM32D_WE_O, n41380, n45079, n70, n10004, n45080, 
            n67, n10006, n64, n10008, n58, n10012, n52, n10016, 
            n49, n10018, n43, n10022, n45076, n40, n10024, n37, 
            n10026, n34, n10028, \selected_1__N_354[0] , LM32D_STB_O, 
            \LM32I_ADR_O[9] , n41390, n30986, n47, \LM32I_ADR_O[14] , 
            \SHAREDBUS_ADR_I[15] , n41234, n61, bus_error_f_N_1884, 
            n41429, \next_cycle_type[2] , n13990, n30900, n41410, 
            REF_CLK_c_enable_97, \LM32I_ADR_O[11] , n41310, n32728, 
            \LM32I_ADR_O[13] , ROM_DAT_O, n8, n8_adj_273, n8_adj_274, 
            n8_adj_275, n8_adj_276, n3, n3_adj_277, n8_adj_278, n3_adj_279, 
            n8_adj_280, n8_adj_281, n3_adj_282, n8_adj_283, n8_adj_284, 
            n8_adj_285, n8_adj_286, n8_adj_287, n3_adj_288, n41255, 
            n15, n35788, n3_adj_289, n3_adj_290, n8_adj_291, n8_adj_292, 
            n8_adj_293, n8_adj_294, LM32D_DAT_O, n41324, data, n69, 
            ebrEBR_DAT_O, \genblk1.write_data_7__N_3573 , n8_adj_296, 
            n8_adj_297, n8_adj_298, n8_adj_299, n8_adj_300, n11, n8_adj_301, 
            n3_adj_302, \LM32I_ADR_O[8] , inst3_Empty, n35204, \reg_04[29] , 
            n33332, \reg_04[4] , n33294, \reg_04[14] , n33370, \reg_04[17] , 
            n33256, \reg_04[22] , n33218, \reg_04[24] , n33180, n41262, 
            n19822, \counter[2] , n8_adj_303, n41344, n41345, n30231, 
            write_enable, \state_1__N_3407[1] , n6362, n41309, n87, 
            \genblk1.write_data_23__N_3541 , \LM32I_ADR_O[6] , \SHAREDBUS_ADR_I[5] , 
            n41275, \LM32I_ADR_O[4] , \SHAREDBUS_ADR_I[29] , n32174, 
            \SHAREDBUS_ADR_I[25] , n35605, \SHAREDBUS_ADR_I[20] , n41289, 
            selected, REF_CLK_c, REF_CLK_c_enable_1606, \LM32D_ADR_O[10] , 
            n46, n41306, \SHAREDBUS_DAT_I[14] , n78, \SHAREDBUS_DAT_I[15] , 
            \SHAREDBUS_DAT_I[10] , \SHAREDBUS_DAT_I[9] , \SHAREDBUS_DAT_I[8] , 
            \SHAREDBUS_DAT_I[12] , \SHAREDBUS_DAT_I[11] , n45101, \SHAREDBUS_DAT_I[13] , 
            LM32D_CYC_O, n41326, locked_N_493, REF_CLK_c_enable_1221, 
            \genblk1.write_data_15__N_3557 , n41292, n41488, LM32D_SEL_O, 
            n41307, n41485, write_ack, n41278, n41328, \SHAREDBUS_DAT_I[31] , 
            \SHAREDBUS_DAT_I[30] , \SHAREDBUS_DAT_I[24] , \SHAREDBUS_DAT_I[28] , 
            \SHAREDBUS_DAT_I[29] , \LM32D_ADR_O[29] , \LM32I_ADR_O[29] , 
            \LM32D_ADR_O[18] , \LM32I_ADR_O[18] , \SHAREDBUS_ADR_I[18] , 
            \LM32D_ADR_O[31] , \LM32I_ADR_O[31] , \SHAREDBUS_ADR_I[31] , 
            \LM32D_ADR_O[27] , \LM32I_ADR_O[27] , \SHAREDBUS_ADR_I[27] , 
            \LM32D_ADR_O[23] , \LM32I_ADR_O[23] , \SHAREDBUS_ADR_I[23] , 
            \LM32I_ADR_O[10] , \SHAREDBUS_ADR_I[10] , n954, \LM32D_ADR_O[15] , 
            \LM32I_ADR_O[15] , \LM32D_ADR_O[26] , \LM32I_ADR_O[26] , \SHAREDBUS_ADR_I[26] , 
            \LM32D_ADR_O[16] , \LM32I_ADR_O[16] , \SHAREDBUS_ADR_I[16] , 
            \LM32D_ADR_O[7] , \LM32I_ADR_O[7] , \SHAREDBUS_ADR_I[7] , 
            \LM32D_ADR_O[25] , \LM32I_ADR_O[25] , n953, \LM32D_ADR_O[5] , 
            \LM32I_ADR_O[5] , \LM32D_ADR_O[20] , \LM32I_ADR_O[20] , \LM32D_ADR_O[24] , 
            \LM32I_ADR_O[24] , \SHAREDBUS_ADR_I[24] , \LM32D_ADR_O[22] , 
            \LM32I_ADR_O[22] , \SHAREDBUS_ADR_I[22] , \LM32D_ADR_O[30] , 
            \LM32I_ADR_O[30] , \SHAREDBUS_ADR_I[30] , \SHAREDBUS_DAT_I[26] , 
            \SHAREDBUS_DAT_I[27] , \SHAREDBUS_DAT_I[25] , write_ack_adj_304, 
            n41243, REF_CLK_c_enable_1581, \LM32D_CTI_O[0] , \LM32I_CTI_O[0] , 
            REF_CLK_c_enable_1597, REF_CLK_c_enable_1605, REF_CLK_c_enable_1589, 
            n41329, n41387, n9, n12390, \LM32D_ADR_O[0] , n71_adj_305, 
            \LM32D_ADR_O[6] , \LM32D_ADR_O[12] , n41346, \LM32I_ADR_O[12] , 
            n41303, \LM32D_ADR_O[4] , \LM32D_ADR_O[9] , n41347, n41222, 
            n41304, n6034, n41330, n41331, n41332, n41333, n41334, 
            n41335, n41336, n41337, n41338, n41339, n41193, REF_CLK_c_enable_1558, 
            n41340, n41341, n41342, n41343, n96, n55, n41279, 
            n29830, REF_CLK_c_enable_1574, \genblk1.write_data_31__N_3525 , 
            n41482, \LM32I_ADR_O[2] , n32216, n61_adj_306, n21, n33, 
            n31955, n32220, n41210, n15_adj_307, n35868, n41225, 
            n19, n41226, n41260, n34816, n11831, n41323, n41239, 
            n41238, REF_CLK_c_enable_1131, n41221, \LM32D_ADR_O[14] , 
            n41298, REF_CLK_c_enable_1550, REF_CLK_c_enable_1566, \LM32D_ADR_O[2] , 
            \LM32D_ADR_O[13] , n41300, \next_cycle_type[2]_adj_308 , \LM32D_ADR_O[11] , 
            n37905, n41299, n37904, \LM32D_ADR_O[8] , n37906, n41301, 
            n37903) /* synthesis syn_module_defined=1 */ ;
    input LM32D_WE_O;
    output n41380;
    output n45079;
    input n70;
    output n10004;
    output n45080;
    input n67;
    output n10006;
    input n64;
    output n10008;
    input n58;
    output n10012;
    input n52;
    output n10016;
    input n49;
    output n10018;
    input n43;
    output n10022;
    output n45076;
    input n40;
    output n10024;
    input n37;
    output n10026;
    input n34;
    output n10028;
    input \selected_1__N_354[0] ;
    input LM32D_STB_O;
    input \LM32I_ADR_O[9] ;
    output n41390;
    input n30986;
    output n47;
    input \LM32I_ADR_O[14] ;
    output \SHAREDBUS_ADR_I[15] ;
    output n41234;
    output n61;
    input bus_error_f_N_1884;
    output n41429;
    input \next_cycle_type[2] ;
    input n13990;
    output n30900;
    input n41410;
    output REF_CLK_c_enable_97;
    input \LM32I_ADR_O[11] ;
    output n41310;
    output n32728;
    input \LM32I_ADR_O[13] ;
    input [31:0]ROM_DAT_O;
    output n8;
    output n8_adj_273;
    output n8_adj_274;
    output n8_adj_275;
    output n8_adj_276;
    output n3;
    output n3_adj_277;
    output n8_adj_278;
    output n3_adj_279;
    output n8_adj_280;
    output n8_adj_281;
    output n3_adj_282;
    output n8_adj_283;
    output n8_adj_284;
    output n8_adj_285;
    output n8_adj_286;
    output n8_adj_287;
    output n3_adj_288;
    output n41255;
    output n15;
    output n35788;
    output n3_adj_289;
    output n3_adj_290;
    output n8_adj_291;
    output n8_adj_292;
    output n8_adj_293;
    output n8_adj_294;
    input [31:0]LM32D_DAT_O;
    output n41324;
    input [31:0]data;
    output [7:0]n69;
    input [31:0]ebrEBR_DAT_O;
    output [7:0]\genblk1.write_data_7__N_3573 ;
    output n8_adj_296;
    output n8_adj_297;
    output n8_adj_298;
    output n8_adj_299;
    output n8_adj_300;
    output n11;
    output n8_adj_301;
    output n3_adj_302;
    input \LM32I_ADR_O[8] ;
    input inst3_Empty;
    output n35204;
    input \reg_04[29] ;
    output n33332;
    input \reg_04[4] ;
    output n33294;
    input \reg_04[14] ;
    output n33370;
    input \reg_04[17] ;
    output n33256;
    input \reg_04[22] ;
    output n33218;
    input \reg_04[24] ;
    output n33180;
    output n41262;
    input n19822;
    input \counter[2] ;
    output n8_adj_303;
    output n41344;
    output n41345;
    output n30231;
    input write_enable;
    input \state_1__N_3407[1] ;
    output n6362;
    output n41309;
    output [7:0]n87;
    output [7:0]\genblk1.write_data_23__N_3541 ;
    input \LM32I_ADR_O[6] ;
    output \SHAREDBUS_ADR_I[5] ;
    output n41275;
    input \LM32I_ADR_O[4] ;
    output \SHAREDBUS_ADR_I[29] ;
    output n32174;
    output \SHAREDBUS_ADR_I[25] ;
    output n35605;
    output \SHAREDBUS_ADR_I[20] ;
    output n41289;
    output [1:0]selected;
    input REF_CLK_c;
    input REF_CLK_c_enable_1606;
    input \LM32D_ADR_O[10] ;
    input n46;
    output n41306;
    output \SHAREDBUS_DAT_I[14] ;
    output [7:0]n78;
    output \SHAREDBUS_DAT_I[15] ;
    output \SHAREDBUS_DAT_I[10] ;
    output \SHAREDBUS_DAT_I[9] ;
    output \SHAREDBUS_DAT_I[8] ;
    output \SHAREDBUS_DAT_I[12] ;
    output \SHAREDBUS_DAT_I[11] ;
    output n45101;
    output \SHAREDBUS_DAT_I[13] ;
    input LM32D_CYC_O;
    output n41326;
    input locked_N_493;
    output REF_CLK_c_enable_1221;
    output [7:0]\genblk1.write_data_15__N_3557 ;
    output n41292;
    output n41488;
    input [3:0]LM32D_SEL_O;
    output n41307;
    output n41485;
    input write_ack;
    output n41278;
    output n41328;
    output \SHAREDBUS_DAT_I[31] ;
    output \SHAREDBUS_DAT_I[30] ;
    output \SHAREDBUS_DAT_I[24] ;
    output \SHAREDBUS_DAT_I[28] ;
    output \SHAREDBUS_DAT_I[29] ;
    input \LM32D_ADR_O[29] ;
    input \LM32I_ADR_O[29] ;
    input \LM32D_ADR_O[18] ;
    input \LM32I_ADR_O[18] ;
    output \SHAREDBUS_ADR_I[18] ;
    input \LM32D_ADR_O[31] ;
    input \LM32I_ADR_O[31] ;
    output \SHAREDBUS_ADR_I[31] ;
    input \LM32D_ADR_O[27] ;
    input \LM32I_ADR_O[27] ;
    output \SHAREDBUS_ADR_I[27] ;
    input \LM32D_ADR_O[23] ;
    input \LM32I_ADR_O[23] ;
    output \SHAREDBUS_ADR_I[23] ;
    input \LM32I_ADR_O[10] ;
    output \SHAREDBUS_ADR_I[10] ;
    output [0:0]n954;
    input \LM32D_ADR_O[15] ;
    input \LM32I_ADR_O[15] ;
    input \LM32D_ADR_O[26] ;
    input \LM32I_ADR_O[26] ;
    output \SHAREDBUS_ADR_I[26] ;
    input \LM32D_ADR_O[16] ;
    input \LM32I_ADR_O[16] ;
    output \SHAREDBUS_ADR_I[16] ;
    input \LM32D_ADR_O[7] ;
    input \LM32I_ADR_O[7] ;
    output \SHAREDBUS_ADR_I[7] ;
    input \LM32D_ADR_O[25] ;
    input \LM32I_ADR_O[25] ;
    output [0:0]n953;
    input \LM32D_ADR_O[5] ;
    input \LM32I_ADR_O[5] ;
    input \LM32D_ADR_O[20] ;
    input \LM32I_ADR_O[20] ;
    input \LM32D_ADR_O[24] ;
    input \LM32I_ADR_O[24] ;
    output \SHAREDBUS_ADR_I[24] ;
    input \LM32D_ADR_O[22] ;
    input \LM32I_ADR_O[22] ;
    output \SHAREDBUS_ADR_I[22] ;
    input \LM32D_ADR_O[30] ;
    input \LM32I_ADR_O[30] ;
    output \SHAREDBUS_ADR_I[30] ;
    output \SHAREDBUS_DAT_I[26] ;
    output \SHAREDBUS_DAT_I[27] ;
    output \SHAREDBUS_DAT_I[25] ;
    input write_ack_adj_304;
    output n41243;
    output REF_CLK_c_enable_1581;
    input \LM32D_CTI_O[0] ;
    input \LM32I_CTI_O[0] ;
    output REF_CLK_c_enable_1597;
    output REF_CLK_c_enable_1605;
    output REF_CLK_c_enable_1589;
    output n41329;
    input n41387;
    output n9;
    output n12390;
    input \LM32D_ADR_O[0] ;
    output n71_adj_305;
    input \LM32D_ADR_O[6] ;
    input \LM32D_ADR_O[12] ;
    output n41346;
    input \LM32I_ADR_O[12] ;
    output n41303;
    input \LM32D_ADR_O[4] ;
    input \LM32D_ADR_O[9] ;
    output n41347;
    output n41222;
    output n41304;
    output n6034;
    output n41330;
    output n41331;
    output n41332;
    output n41333;
    output n41334;
    output n41335;
    output n41336;
    output n41337;
    output n41338;
    output n41339;
    input n41193;
    output REF_CLK_c_enable_1558;
    output n41340;
    output n41341;
    output n41342;
    output n41343;
    output [7:0]n96;
    input n55;
    input n41279;
    output n29830;
    output REF_CLK_c_enable_1574;
    output [7:0]\genblk1.write_data_31__N_3525 ;
    output n41482;
    input \LM32I_ADR_O[2] ;
    output n32216;
    input n61_adj_306;
    input n21;
    output n33;
    input n31955;
    output n32220;
    input n41210;
    input n15_adj_307;
    input n35868;
    input n41225;
    input n19;
    input n41226;
    input n41260;
    input n34816;
    output n11831;
    output n41323;
    output n41239;
    output n41238;
    output REF_CLK_c_enable_1131;
    output n41221;
    input \LM32D_ADR_O[14] ;
    output n41298;
    output REF_CLK_c_enable_1550;
    output REF_CLK_c_enable_1566;
    input \LM32D_ADR_O[2] ;
    input \LM32D_ADR_O[13] ;
    output n41300;
    input \next_cycle_type[2]_adj_308 ;
    input \LM32D_ADR_O[11] ;
    output n37905;
    output n41299;
    output n37904;
    input \LM32D_ADR_O[8] ;
    output n37906;
    output n41301;
    output n37903;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    
    wire n45082, n45081, n45074, n45077, n45073, n45072, n45071, 
        n41386, n9234, REF_CLK_c_enable_1237, n41427, n41256, REF_CLK_c_enable_1623, 
        n36341, n41481;
    wire [1:0]selected_1__N_350;
    
    wire n45097, n41480, n41486, n41487, n41483, n41484, n18080, 
        n45084, n45083, n38693, n34850, n34836;
    
    LUT4 i4672_3_lut_4_lut (.A(LM32D_WE_O), .B(n41380), .C(n45079), .D(n70), 
         .Z(n10004)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i4672_3_lut_4_lut.init = 16'hf780;
    LUT4 i4674_3_lut_4_lut (.A(LM32D_WE_O), .B(n41380), .C(n45080), .D(n67), 
         .Z(n10006)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i4674_3_lut_4_lut.init = 16'hf780;
    LUT4 i4676_3_lut_4_lut (.A(LM32D_WE_O), .B(n41380), .C(n45082), .D(n64), 
         .Z(n10008)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i4676_3_lut_4_lut.init = 16'hf780;
    LUT4 i4680_3_lut_4_lut (.A(LM32D_WE_O), .B(n41380), .C(n45081), .D(n58), 
         .Z(n10012)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i4680_3_lut_4_lut.init = 16'hf780;
    LUT4 i4684_3_lut_4_lut (.A(LM32D_WE_O), .B(n41380), .C(n45074), .D(n52), 
         .Z(n10016)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i4684_3_lut_4_lut.init = 16'hf780;
    LUT4 i4686_3_lut_4_lut (.A(LM32D_WE_O), .B(n41380), .C(n45077), .D(n49), 
         .Z(n10018)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i4686_3_lut_4_lut.init = 16'hf780;
    LUT4 i4690_3_lut_4_lut (.A(LM32D_WE_O), .B(n41380), .C(n45073), .D(n43), 
         .Z(n10022)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i4690_3_lut_4_lut.init = 16'hf780;
    LUT4 i6_3_lut_4_lut (.A(LM32D_WE_O), .B(n41380), .C(n45076), .D(n40), 
         .Z(n10024)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i6_3_lut_4_lut.init = 16'hf780;
    LUT4 i4694_3_lut_4_lut (.A(LM32D_WE_O), .B(n41380), .C(n45072), .D(n37), 
         .Z(n10026)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i4694_3_lut_4_lut.init = 16'hf780;
    LUT4 i4696_3_lut_4_lut (.A(LM32D_WE_O), .B(n41380), .C(n45071), .D(n34), 
         .Z(n10028)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i4696_3_lut_4_lut.init = 16'hf780;
    LUT4 i33072_3_lut_4_lut (.A(\selected_1__N_354[0] ), .B(n41386), .C(LM32D_STB_O), 
         .D(n9234), .Z(REF_CLK_c_enable_1237)) /* synthesis lut_function=(A ((D)+!B)+!A (B (D)+!B (C))) */ ;
    defparam i33072_3_lut_4_lut.init = 16'hfe32;
    LUT4 i1_2_lut_4_lut (.A(\LM32I_ADR_O[9] ), .B(n45077), .C(n41390), 
         .D(n30986), .Z(n47)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_4_lut.init = 16'hff35;
    LUT4 i1_2_lut_rep_829_4_lut (.A(\LM32I_ADR_O[14] ), .B(n45071), .C(n41390), 
         .D(\SHAREDBUS_ADR_I[15] ), .Z(n41234)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_rep_829_4_lut.init = 16'hffca;
    LUT4 i1_2_lut_4_lut_adj_654 (.A(\LM32I_ADR_O[14] ), .B(n45071), .C(n41390), 
         .D(\SHAREDBUS_ADR_I[15] ), .Z(n61)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_4_lut_adj_654.init = 16'hff35;
    LUT4 i1_3_lut_4_lut (.A(bus_error_f_N_1884), .B(n41429), .C(\next_cycle_type[2] ), 
         .D(n13990), .Z(n30900)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam i1_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(bus_error_f_N_1884), .B(n41429), 
         .C(n13990), .D(n41410), .Z(REF_CLK_c_enable_97)) /* synthesis lut_function=(A (B (C))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'hd580;
    LUT4 i1_2_lut_4_lut_adj_655 (.A(\LM32I_ADR_O[11] ), .B(n45073), .C(n41390), 
         .D(n41310), .Z(n32728)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_4_lut_adj_655.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut (.A(\LM32I_ADR_O[13] ), .B(n45072), .C(n41390), 
         .D(ROM_DAT_O[4]), .Z(n8)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_656 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[29]), .Z(n8_adj_273)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_656.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_657 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[30]), .Z(n8_adj_274)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_657.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_658 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[8]), .Z(n8_adj_275)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_658.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_659 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[26]), .Z(n8_adj_276)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_659.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_660 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[9]), .Z(n3)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_660.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_661 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[13]), .Z(n3_adj_277)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_661.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_662 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[12]), .Z(n8_adj_278)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_662.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_663 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[11]), .Z(n3_adj_279)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_663.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_664 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[1]), .Z(n8_adj_280)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_664.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_665 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[19]), .Z(n8_adj_281)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_665.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_666 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[18]), .Z(n3_adj_282)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_666.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_667 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[2]), .Z(n8_adj_283)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_667.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_668 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[3]), .Z(n8_adj_284)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_668.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_669 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[0]), .Z(n8_adj_285)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_669.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_670 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[31]), .Z(n8_adj_286)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_670.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_671 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[17]), .Z(n8_adj_287)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_671.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_672 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[25]), .Z(n3_adj_288)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_672.init = 16'h3500;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n41427), .B(n41390), .C(n41256), .D(n41255), 
         .Z(n15)) /* synthesis lut_function=(A (B (C+!(D))+!B (C+(D)))+!A (C+(D))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf7f8;
    LUT4 i30626_2_lut_3_lut_4_lut (.A(n41427), .B(n41390), .C(n41256), 
         .D(n41255), .Z(n35788)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C+(D))) */ ;
    defparam i30626_2_lut_3_lut_4_lut.init = 16'hf7f0;
    LUT4 i1_2_lut_2_lut_4_lut_adj_673 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[21]), .Z(n3_adj_289)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_673.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_674 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[28]), .Z(n3_adj_290)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_674.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_675 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[6]), .Z(n8_adj_291)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_675.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_676 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[22]), .Z(n8_adj_292)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_676.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_677 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[7]), .Z(n8_adj_293)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_677.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_678 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[10]), .Z(n8_adj_294)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_678.init = 16'h3500;
    LUT4 mux_6_i1_3_lut_4_lut (.A(LM32D_DAT_O[0]), .B(n41380), .C(n41324), 
         .D(data[0]), .Z(n69[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam mux_6_i1_3_lut_4_lut.init = 16'h8f80;
    LUT4 EBR_DAT_O_7__I_0_i1_3_lut_4_lut (.A(LM32D_DAT_O[0]), .B(n41380), 
         .C(n41324), .D(ebrEBR_DAT_O[0]), .Z(\genblk1.write_data_7__N_3573 [0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam EBR_DAT_O_7__I_0_i1_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_2_lut_4_lut_adj_679 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[23]), .Z(n8_adj_296)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_679.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_680 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[5]), .Z(n8_adj_297)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_680.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_681 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[16]), .Z(n8_adj_298)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_681.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_682 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[20]), .Z(n8_adj_299)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_682.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_683 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[27]), .Z(n8_adj_300)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_683.init = 16'h3500;
    LUT4 i1_2_lut_2_lut_4_lut_adj_684 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[24]), .Z(n11)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_684.init = 16'h3500;
    LUT4 mux_6_i2_3_lut_4_lut (.A(LM32D_DAT_O[1]), .B(n41380), .C(n41324), 
         .D(data[1]), .Z(n69[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam mux_6_i2_3_lut_4_lut.init = 16'h8f80;
    LUT4 EBR_DAT_O_7__I_0_i2_3_lut_4_lut (.A(LM32D_DAT_O[1]), .B(n41380), 
         .C(n41324), .D(ebrEBR_DAT_O[1]), .Z(\genblk1.write_data_7__N_3573 [1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam EBR_DAT_O_7__I_0_i2_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_6_i3_3_lut_4_lut (.A(LM32D_DAT_O[2]), .B(n41380), .C(n41324), 
         .D(data[2]), .Z(n69[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam mux_6_i3_3_lut_4_lut.init = 16'h8f80;
    LUT4 EBR_DAT_O_7__I_0_i3_3_lut_4_lut (.A(LM32D_DAT_O[2]), .B(n41380), 
         .C(n41324), .D(ebrEBR_DAT_O[2]), .Z(\genblk1.write_data_7__N_3573 [2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam EBR_DAT_O_7__I_0_i3_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_2_lut_4_lut_adj_685 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[14]), .Z(n8_adj_301)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_685.init = 16'h3500;
    LUT4 mux_6_i4_3_lut_4_lut (.A(LM32D_DAT_O[3]), .B(n41380), .C(n41324), 
         .D(data[3]), .Z(n69[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam mux_6_i4_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_2_lut_4_lut_adj_686 (.A(\LM32I_ADR_O[13] ), .B(n45072), 
         .C(n41390), .D(ROM_DAT_O[15]), .Z(n3_adj_302)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_2_lut_4_lut_adj_686.init = 16'h3500;
    LUT4 i1_2_lut_4_lut_adj_687 (.A(\LM32I_ADR_O[8] ), .B(n45074), .C(n41390), 
         .D(inst3_Empty), .Z(n35204)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_4_lut_adj_687.init = 16'h00ca;
    LUT4 i1_2_lut_4_lut_adj_688 (.A(\LM32I_ADR_O[8] ), .B(n45074), .C(n41390), 
         .D(\reg_04[29] ), .Z(n33332)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_4_lut_adj_688.init = 16'hca00;
    LUT4 EBR_DAT_O_7__I_0_i4_3_lut_4_lut (.A(LM32D_DAT_O[3]), .B(n41380), 
         .C(n41324), .D(ebrEBR_DAT_O[3]), .Z(\genblk1.write_data_7__N_3573 [3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam EBR_DAT_O_7__I_0_i4_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13767_3_lut_4_lut (.A(LM32D_DAT_O[4]), .B(n41380), .C(n41324), 
         .D(ebrEBR_DAT_O[4]), .Z(\genblk1.write_data_7__N_3573 [4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam i13767_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_4_lut_adj_689 (.A(\LM32I_ADR_O[8] ), .B(n45074), .C(n41390), 
         .D(\reg_04[4] ), .Z(n33294)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_4_lut_adj_689.init = 16'hca00;
    LUT4 i1_2_lut_4_lut_adj_690 (.A(\LM32I_ADR_O[8] ), .B(n45074), .C(n41390), 
         .D(\reg_04[14] ), .Z(n33370)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_4_lut_adj_690.init = 16'hca00;
    LUT4 i1_2_lut_4_lut_adj_691 (.A(\LM32I_ADR_O[8] ), .B(n45074), .C(n41390), 
         .D(\reg_04[17] ), .Z(n33256)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_4_lut_adj_691.init = 16'hca00;
    LUT4 i1_2_lut_4_lut_adj_692 (.A(\LM32I_ADR_O[8] ), .B(n45074), .C(n41390), 
         .D(\reg_04[22] ), .Z(n33218)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_4_lut_adj_692.init = 16'hca00;
    LUT4 i1_2_lut_4_lut_adj_693 (.A(\LM32I_ADR_O[8] ), .B(n45074), .C(n41390), 
         .D(\reg_04[24] ), .Z(n33180)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_4_lut_adj_693.init = 16'hca00;
    LUT4 i1_2_lut_rep_857_4_lut (.A(\LM32I_ADR_O[8] ), .B(n45074), .C(n41390), 
         .D(n41310), .Z(n41262)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_rep_857_4_lut.init = 16'hca00;
    LUT4 mux_6_i5_3_lut_4_lut (.A(LM32D_DAT_O[4]), .B(n41380), .C(n41324), 
         .D(data[4]), .Z(n69[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam mux_6_i5_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_6_i6_3_lut_4_lut (.A(LM32D_DAT_O[5]), .B(n41380), .C(n41324), 
         .D(data[5]), .Z(n69[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam mux_6_i6_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_3_lut_4_lut_adj_694 (.A(LM32D_WE_O), .B(n41380), .C(n19822), 
         .D(\counter[2] ), .Z(n8_adj_303)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i1_2_lut_3_lut_4_lut_adj_694.init = 16'h7000;
    LUT4 i33152_2_lut_3_lut_4_lut (.A(LM32D_WE_O), .B(n41380), .C(n41344), 
         .D(n41345), .Z(n30231)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i33152_2_lut_3_lut_4_lut.init = 16'h0007;
    LUT4 EBR_DAT_O_7__I_0_i6_3_lut_4_lut (.A(LM32D_DAT_O[5]), .B(n41380), 
         .C(n41324), .D(ebrEBR_DAT_O[5]), .Z(\genblk1.write_data_7__N_3573 [5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam EBR_DAT_O_7__I_0_i6_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_3_lut_4_lut_adj_695 (.A(LM32D_WE_O), .B(n41380), .C(write_enable), 
         .D(\state_1__N_3407[1] ), .Z(n6362)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i1_3_lut_4_lut_adj_695.init = 16'hf800;
    LUT4 mux_6_i7_3_lut_4_lut (.A(LM32D_DAT_O[6]), .B(n41380), .C(n41324), 
         .D(data[6]), .Z(n69[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam mux_6_i7_3_lut_4_lut.init = 16'h8f80;
    LUT4 EBR_DAT_O_7__I_0_i7_3_lut_4_lut (.A(LM32D_DAT_O[6]), .B(n41380), 
         .C(n41324), .D(ebrEBR_DAT_O[6]), .Z(\genblk1.write_data_7__N_3573 [6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam EBR_DAT_O_7__I_0_i7_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_6_i8_3_lut_4_lut (.A(LM32D_DAT_O[7]), .B(n41380), .C(n41324), 
         .D(data[7]), .Z(n69[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam mux_6_i8_3_lut_4_lut.init = 16'h8f80;
    LUT4 EBR_DAT_O_7__I_0_i8_3_lut_4_lut (.A(LM32D_DAT_O[7]), .B(n41380), 
         .C(n41324), .D(ebrEBR_DAT_O[7]), .Z(\genblk1.write_data_7__N_3573 [7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam EBR_DAT_O_7__I_0_i8_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_8_i1_3_lut_4_lut (.A(LM32D_DAT_O[16]), .B(n41380), .C(n41309), 
         .D(data[16]), .Z(n87[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam mux_8_i1_3_lut_4_lut.init = 16'h8f80;
    LUT4 EBR_DAT_O_23__I_0_i1_3_lut_4_lut (.A(LM32D_DAT_O[16]), .B(n41380), 
         .C(n41309), .D(ebrEBR_DAT_O[16]), .Z(\genblk1.write_data_23__N_3541 [0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam EBR_DAT_O_23__I_0_i1_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_8_i2_3_lut_4_lut (.A(LM32D_DAT_O[17]), .B(n41380), .C(n41309), 
         .D(data[17]), .Z(n87[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam mux_8_i2_3_lut_4_lut.init = 16'h8f80;
    LUT4 EBR_DAT_O_23__I_0_i2_3_lut_4_lut (.A(LM32D_DAT_O[17]), .B(n41380), 
         .C(n41309), .D(ebrEBR_DAT_O[17]), .Z(\genblk1.write_data_23__N_3541 [1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam EBR_DAT_O_23__I_0_i2_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_8_i3_3_lut_4_lut (.A(LM32D_DAT_O[18]), .B(n41380), .C(n41309), 
         .D(data[18]), .Z(n87[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam mux_8_i3_3_lut_4_lut.init = 16'h8f80;
    LUT4 EBR_DAT_O_23__I_0_i3_3_lut_4_lut (.A(LM32D_DAT_O[18]), .B(n41380), 
         .C(n41309), .D(ebrEBR_DAT_O[18]), .Z(\genblk1.write_data_23__N_3541 [2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam EBR_DAT_O_23__I_0_i3_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_8_i4_3_lut_4_lut (.A(LM32D_DAT_O[19]), .B(n41380), .C(n41309), 
         .D(data[19]), .Z(n87[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam mux_8_i4_3_lut_4_lut.init = 16'h8f80;
    LUT4 EBR_DAT_O_23__I_0_i4_3_lut_4_lut (.A(LM32D_DAT_O[19]), .B(n41380), 
         .C(n41309), .D(ebrEBR_DAT_O[19]), .Z(\genblk1.write_data_23__N_3541 [3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam EBR_DAT_O_23__I_0_i4_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13240_3_lut_4_lut (.A(LM32D_DAT_O[20]), .B(n41380), .C(n41309), 
         .D(ebrEBR_DAT_O[20]), .Z(\genblk1.write_data_23__N_3541 [4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam i13240_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_8_i5_3_lut_4_lut (.A(LM32D_DAT_O[20]), .B(n41380), .C(n41309), 
         .D(data[20]), .Z(n87[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam mux_8_i5_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_8_i6_3_lut_4_lut (.A(LM32D_DAT_O[21]), .B(n41380), .C(n41309), 
         .D(data[21]), .Z(n87[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam mux_8_i6_3_lut_4_lut.init = 16'h8f80;
    LUT4 EBR_DAT_O_23__I_0_i6_3_lut_4_lut (.A(LM32D_DAT_O[21]), .B(n41380), 
         .C(n41309), .D(ebrEBR_DAT_O[21]), .Z(\genblk1.write_data_23__N_3541 [5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam EBR_DAT_O_23__I_0_i6_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_8_i7_3_lut_4_lut (.A(LM32D_DAT_O[22]), .B(n41380), .C(n41309), 
         .D(data[22]), .Z(n87[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam mux_8_i7_3_lut_4_lut.init = 16'h8f80;
    LUT4 EBR_DAT_O_23__I_0_i7_3_lut_4_lut (.A(LM32D_DAT_O[22]), .B(n41380), 
         .C(n41309), .D(ebrEBR_DAT_O[22]), .Z(\genblk1.write_data_23__N_3541 [6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam EBR_DAT_O_23__I_0_i7_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_8_i8_3_lut_4_lut (.A(LM32D_DAT_O[23]), .B(n41380), .C(n41309), 
         .D(data[23]), .Z(n87[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam mux_8_i8_3_lut_4_lut.init = 16'h8f80;
    LUT4 EBR_DAT_O_23__I_0_i8_3_lut_4_lut (.A(LM32D_DAT_O[23]), .B(n41380), 
         .C(n41309), .D(ebrEBR_DAT_O[23]), .Z(\genblk1.write_data_23__N_3541 [7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(284[2] 285[4])
    defparam EBR_DAT_O_23__I_0_i8_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_rep_870_4_lut (.A(\LM32I_ADR_O[6] ), .B(n45081), .C(n41390), 
         .D(\SHAREDBUS_ADR_I[5] ), .Z(n41275)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_rep_870_4_lut.init = 16'hffca;
    LUT4 i1_2_lut_4_lut_adj_696 (.A(\LM32I_ADR_O[4] ), .B(n45082), .C(n41390), 
         .D(\SHAREDBUS_ADR_I[29] ), .Z(n32174)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_4_lut_adj_696.init = 16'hffca;
    LUT4 i30460_2_lut_4_lut (.A(\LM32I_ADR_O[4] ), .B(n45082), .C(n41390), 
         .D(\SHAREDBUS_ADR_I[25] ), .Z(n35605)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i30460_2_lut_4_lut.init = 16'hffca;
    LUT4 i1_2_lut_rep_884_4_lut (.A(\LM32I_ADR_O[4] ), .B(n45082), .C(n41390), 
         .D(\SHAREDBUS_ADR_I[20] ), .Z(n41289)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(279[2] 281[5])
    defparam i1_2_lut_rep_884_4_lut.init = 16'hffca;
    FD1P3DX selected_i1 (.D(n36341), .SP(REF_CLK_c_enable_1623), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(selected[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=1, LSE_RCOL=20, LSE_LLINE=488, LSE_RLINE=529 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(252[7] 275[5])
    defparam selected_i1.GSR = "ENABLED";
    LUT4 i4688_3_lut_4_lut_then_4_lut (.A(\LM32D_ADR_O[10] ), .B(selected[0]), 
         .C(selected[1]), .D(n46), .Z(n41481)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (B (D)+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i4688_3_lut_4_lut_then_4_lut.init = 16'hef20;
    FD1P3DX selected_i0_rep_1063 (.D(selected_1__N_350[0]), .SP(REF_CLK_c_enable_1237), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(n45097)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=1, LSE_RCOL=20, LSE_LLINE=488, LSE_RLINE=529 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(252[7] 275[5])
    defparam selected_i0_rep_1063.GSR = "ENABLED";
    LUT4 i4688_3_lut_4_lut_else_4_lut (.A(n46), .Z(n41480)) /* synthesis lut_function=(A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i4688_3_lut_4_lut_else_4_lut.init = 16'haaaa;
    LUT4 mux_7_i7_3_lut_4_lut (.A(n41429), .B(n41306), .C(\SHAREDBUS_DAT_I[14] ), 
         .D(data[14]), .Z(n78[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_7_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_7_i8_3_lut_4_lut (.A(n41429), .B(n41306), .C(\SHAREDBUS_DAT_I[15] ), 
         .D(data[15]), .Z(n78[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_7_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_7_i3_3_lut_4_lut (.A(n41429), .B(n41306), .C(\SHAREDBUS_DAT_I[10] ), 
         .D(data[10]), .Z(n78[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_7_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_7_i2_3_lut_4_lut (.A(n41429), .B(n41306), .C(\SHAREDBUS_DAT_I[9] ), 
         .D(data[9]), .Z(n78[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_7_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_7_i1_3_lut_4_lut (.A(n41429), .B(n41306), .C(\SHAREDBUS_DAT_I[8] ), 
         .D(data[8]), .Z(n78[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_7_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_7_i5_3_lut_4_lut (.A(n41429), .B(n41306), .C(\SHAREDBUS_DAT_I[12] ), 
         .D(data[12]), .Z(n78[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_7_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_7_i4_3_lut_4_lut (.A(n41429), .B(n41306), .C(\SHAREDBUS_DAT_I[11] ), 
         .D(data[11]), .Z(n78[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_7_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_975 (.A(n45097), .B(n45101), .Z(n41380)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_rep_975.init = 16'h4444;
    LUT4 mux_7_i6_3_lut_4_lut (.A(n41429), .B(n41306), .C(\SHAREDBUS_DAT_I[13] ), 
         .D(data[13]), .Z(n78[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_7_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_921_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_CYC_O), 
         .Z(n41326)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_rep_921_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_rep_764_3_lut_4_lut (.A(selected[0]), .B(selected[1]), 
         .C(locked_N_493), .D(LM32D_CYC_O), .Z(REF_CLK_c_enable_1221)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_rep_764_3_lut_4_lut.init = 16'h4000;
    LUT4 EBR_DAT_O_15__I_0_i1_3_lut_4_lut (.A(n41429), .B(n41306), .C(\SHAREDBUS_DAT_I[8] ), 
         .D(ebrEBR_DAT_O[8]), .Z(\genblk1.write_data_15__N_3557 [0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam EBR_DAT_O_15__I_0_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_887_3_lut_4_lut (.A(selected[0]), .B(selected[1]), 
         .C(\counter[2] ), .D(LM32D_WE_O), .Z(n41292)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C))) */ ;
    defparam i1_2_lut_rep_887_3_lut_4_lut.init = 16'hb0f0;
    PFUMX i34377 (.BLUT(n41486), .ALUT(n41487), .C0(LM32D_WE_O), .Z(n41488));
    LUT4 i1_2_lut_rep_901_3_lut (.A(n45097), .B(n45101), .C(LM32D_SEL_O[1]), 
         .Z(n41306)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_rep_901_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_rep_902_3_lut (.A(n45097), .B(n45101), .C(LM32D_SEL_O[3]), 
         .Z(n41307)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_rep_902_3_lut.init = 16'h4040;
    PFUMX i34375 (.BLUT(n41483), .ALUT(n41484), .C0(LM32D_WE_O), .Z(n41485));
    LUT4 EBR_DAT_O_15__I_0_i7_3_lut_4_lut (.A(n41429), .B(n41306), .C(\SHAREDBUS_DAT_I[14] ), 
         .D(ebrEBR_DAT_O[14]), .Z(\genblk1.write_data_15__N_3557 [6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam EBR_DAT_O_15__I_0_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_873_3_lut_4_lut (.A(n45097), .B(n45101), .C(write_ack), 
         .D(LM32D_WE_O), .Z(n41278)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_rep_873_3_lut_4_lut.init = 16'h0400;
    LUT4 i14513_2_lut_rep_923_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[0]), 
         .Z(n41328)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14513_2_lut_rep_923_3_lut.init = 16'h4040;
    LUT4 i14914_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[31]), 
         .Z(\SHAREDBUS_DAT_I[31] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14914_2_lut_3_lut.init = 16'h4040;
    LUT4 i14913_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[30]), 
         .Z(\SHAREDBUS_DAT_I[30] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14913_2_lut_3_lut.init = 16'h4040;
    LUT4 EBR_DAT_O_15__I_0_i6_3_lut_4_lut (.A(n41429), .B(n41306), .C(\SHAREDBUS_DAT_I[13] ), 
         .D(ebrEBR_DAT_O[13]), .Z(\genblk1.write_data_15__N_3557 [5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam EBR_DAT_O_15__I_0_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i14907_2_lut_3_lut (.A(selected[0]), .B(n45101), .C(LM32D_DAT_O[24]), 
         .Z(\SHAREDBUS_DAT_I[24] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14907_2_lut_3_lut.init = 16'h4040;
    LUT4 i14898_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[15]), 
         .Z(\SHAREDBUS_DAT_I[15] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14898_2_lut_3_lut.init = 16'h4040;
    LUT4 i14897_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[14]), 
         .Z(\SHAREDBUS_DAT_I[14] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14897_2_lut_3_lut.init = 16'h4040;
    LUT4 EBR_DAT_O_15__I_0_i5_3_lut_4_lut (.A(n41429), .B(n41306), .C(\SHAREDBUS_DAT_I[12] ), 
         .D(ebrEBR_DAT_O[12]), .Z(\genblk1.write_data_15__N_3557 [4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam EBR_DAT_O_15__I_0_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i14911_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[28]), 
         .Z(\SHAREDBUS_DAT_I[28] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14911_2_lut_3_lut.init = 16'h4040;
    LUT4 i14892_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[9]), 
         .Z(\SHAREDBUS_DAT_I[9] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14892_2_lut_3_lut.init = 16'h4040;
    LUT4 i14894_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[11]), 
         .Z(\SHAREDBUS_DAT_I[11] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14894_2_lut_3_lut.init = 16'h4040;
    LUT4 i14912_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[29]), 
         .Z(\SHAREDBUS_DAT_I[29] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14912_2_lut_3_lut.init = 16'h4040;
    LUT4 i14895_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[12]), 
         .Z(\SHAREDBUS_DAT_I[12] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14895_2_lut_3_lut.init = 16'h4040;
    LUT4 i14893_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[10]), 
         .Z(\SHAREDBUS_DAT_I[10] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14893_2_lut_3_lut.init = 16'h4040;
    LUT4 i14891_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[8]), 
         .Z(\SHAREDBUS_DAT_I[8] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14891_2_lut_3_lut.init = 16'h4040;
    LUT4 WBS_ADR_I_31__I_0_i30_4_lut_4_lut_4_lut (.A(n45097), .B(n45101), 
         .C(\LM32D_ADR_O[29] ), .D(\LM32I_ADR_O[29] ), .Z(\SHAREDBUS_ADR_I[29] )) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam WBS_ADR_I_31__I_0_i30_4_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 WBS_ADR_I_31__I_0_i19_4_lut_4_lut_4_lut (.A(n45097), .B(n45101), 
         .C(\LM32D_ADR_O[18] ), .D(\LM32I_ADR_O[18] ), .Z(\SHAREDBUS_ADR_I[18] )) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam WBS_ADR_I_31__I_0_i19_4_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 WBS_ADR_I_31__I_0_i32_4_lut_4_lut_4_lut (.A(n45097), .B(n45101), 
         .C(\LM32D_ADR_O[31] ), .D(\LM32I_ADR_O[31] ), .Z(\SHAREDBUS_ADR_I[31] )) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam WBS_ADR_I_31__I_0_i32_4_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 WBS_ADR_I_31__I_0_i28_4_lut_4_lut_4_lut (.A(n45097), .B(selected[1]), 
         .C(\LM32D_ADR_O[27] ), .D(\LM32I_ADR_O[27] ), .Z(\SHAREDBUS_ADR_I[27] )) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam WBS_ADR_I_31__I_0_i28_4_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 WBS_ADR_I_31__I_0_i24_4_lut_4_lut_4_lut (.A(selected[0]), .B(selected[1]), 
         .C(\LM32D_ADR_O[23] ), .D(\LM32I_ADR_O[23] ), .Z(\SHAREDBUS_ADR_I[23] )) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam WBS_ADR_I_31__I_0_i24_4_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 WBS_ADR_I_31__I_0_i11_3_lut_4_lut_4_lut (.A(selected[0]), .B(selected[1]), 
         .C(\LM32D_ADR_O[10] ), .D(\LM32I_ADR_O[10] ), .Z(\SHAREDBUS_ADR_I[10] )) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam WBS_ADR_I_31__I_0_i11_3_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 mux_14_i1_4_lut_4_lut_4_lut (.A(selected[0]), .B(n45101), .C(LM32D_STB_O), 
         .D(\selected_1__N_354[0] ), .Z(n954[0])) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_14_i1_4_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 WBS_ADR_I_31__I_0_i16_4_lut_4_lut_4_lut (.A(n45097), .B(n45101), 
         .C(\LM32D_ADR_O[15] ), .D(\LM32I_ADR_O[15] ), .Z(\SHAREDBUS_ADR_I[15] )) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam WBS_ADR_I_31__I_0_i16_4_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 WBS_ADR_I_31__I_0_i27_4_lut_4_lut_4_lut (.A(n45097), .B(n45101), 
         .C(\LM32D_ADR_O[26] ), .D(\LM32I_ADR_O[26] ), .Z(\SHAREDBUS_ADR_I[26] )) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam WBS_ADR_I_31__I_0_i27_4_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 WBS_ADR_I_31__I_0_i17_4_lut_4_lut_4_lut (.A(n45097), .B(n45101), 
         .C(\LM32D_ADR_O[16] ), .D(\LM32I_ADR_O[16] ), .Z(\SHAREDBUS_ADR_I[16] )) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam WBS_ADR_I_31__I_0_i17_4_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 WBS_ADR_I_31__I_0_i8_3_lut_4_lut_4_lut (.A(n45097), .B(n45101), 
         .C(\LM32D_ADR_O[7] ), .D(\LM32I_ADR_O[7] ), .Z(\SHAREDBUS_ADR_I[7] )) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam WBS_ADR_I_31__I_0_i8_3_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 WBS_ADR_I_31__I_0_i26_4_lut_4_lut_4_lut (.A(n45097), .B(n45101), 
         .C(\LM32D_ADR_O[25] ), .D(\LM32I_ADR_O[25] ), .Z(\SHAREDBUS_ADR_I[25] )) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam WBS_ADR_I_31__I_0_i26_4_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 mux_13_i1_4_lut_4_lut_4_lut (.A(n45097), .B(selected[1]), .C(LM32D_CYC_O), 
         .D(bus_error_f_N_1884), .Z(n953[0])) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_13_i1_4_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 WBS_ADR_I_31__I_0_i6_3_lut_4_lut_4_lut (.A(n45097), .B(n45101), 
         .C(\LM32D_ADR_O[5] ), .D(\LM32I_ADR_O[5] ), .Z(\SHAREDBUS_ADR_I[5] )) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam WBS_ADR_I_31__I_0_i6_3_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 WBS_ADR_I_31__I_0_i21_4_lut_4_lut_4_lut (.A(n45097), .B(n45101), 
         .C(\LM32D_ADR_O[20] ), .D(\LM32I_ADR_O[20] ), .Z(\SHAREDBUS_ADR_I[20] )) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam WBS_ADR_I_31__I_0_i21_4_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 WBS_ADR_I_31__I_0_i25_4_lut_4_lut_4_lut (.A(selected[0]), .B(selected[1]), 
         .C(\LM32D_ADR_O[24] ), .D(\LM32I_ADR_O[24] ), .Z(\SHAREDBUS_ADR_I[24] )) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam WBS_ADR_I_31__I_0_i25_4_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 WBS_ADR_I_31__I_0_i23_4_lut_4_lut_4_lut (.A(n45097), .B(n45101), 
         .C(\LM32D_ADR_O[22] ), .D(\LM32I_ADR_O[22] ), .Z(\SHAREDBUS_ADR_I[22] )) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam WBS_ADR_I_31__I_0_i23_4_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 WBS_ADR_I_31__I_0_i31_4_lut_4_lut_4_lut (.A(n45097), .B(n45101), 
         .C(\LM32D_ADR_O[30] ), .D(\LM32I_ADR_O[30] ), .Z(\SHAREDBUS_ADR_I[30] )) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam WBS_ADR_I_31__I_0_i31_4_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 EBR_DAT_O_15__I_0_i4_3_lut_4_lut (.A(n41429), .B(n41306), .C(\SHAREDBUS_DAT_I[11] ), 
         .D(ebrEBR_DAT_O[11]), .Z(\genblk1.write_data_15__N_3557 [3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam EBR_DAT_O_15__I_0_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i14909_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[26]), 
         .Z(\SHAREDBUS_DAT_I[26] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14909_2_lut_3_lut.init = 16'h4040;
    LUT4 EBR_DAT_O_15__I_0_i8_3_lut_4_lut (.A(n41429), .B(n41306), .C(\SHAREDBUS_DAT_I[15] ), 
         .D(ebrEBR_DAT_O[15]), .Z(\genblk1.write_data_15__N_3557 [7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam EBR_DAT_O_15__I_0_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i14910_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[27]), 
         .Z(\SHAREDBUS_DAT_I[27] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14910_2_lut_3_lut.init = 16'h4040;
    LUT4 i14896_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[13]), 
         .Z(\SHAREDBUS_DAT_I[13] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14896_2_lut_3_lut.init = 16'h4040;
    LUT4 i14908_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[25]), 
         .Z(\SHAREDBUS_DAT_I[25] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14908_2_lut_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_rep_838_3_lut_4_lut (.A(n45097), .B(n45101), .C(write_ack_adj_304), 
         .D(LM32D_WE_O), .Z(n41243)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_rep_838_3_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_4_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_SEL_O[0]), 
         .D(n18080), .Z(REF_CLK_c_enable_1581)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C (D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam i1_2_lut_4_lut_4_lut.init = 16'h6200;
    LUT4 i1_4_lut_then_4_lut (.A(locked_N_493), .B(\LM32D_CTI_O[0] ), .C(selected[1]), 
         .D(selected[0]), .Z(n45084)) /* synthesis lut_function=(!((B (C (D)+!C !(D))+!B (C+!(D)))+!A)) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h0a80;
    LUT4 i1_4_lut_else_4_lut (.A(locked_N_493), .B(\LM32D_CTI_O[0] ), .C(selected[1]), 
         .D(selected[0]), .Z(n45083)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h0080;
    LUT4 mux_12_i1_3_lut_rep_850_4_lut_4_lut (.A(\LM32D_CTI_O[0] ), .B(selected[0]), 
         .C(selected[1]), .D(\LM32I_CTI_O[0] ), .Z(n41255)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(296[2] 297[4])
    defparam mux_12_i1_3_lut_rep_850_4_lut_4_lut.init = 16'h2c20;
    FD1P3DX selected_i0 (.D(selected_1__N_350[0]), .SP(REF_CLK_c_enable_1237), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(selected[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=1, LSE_RCOL=20, LSE_LLINE=488, LSE_RLINE=529 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(252[7] 275[5])
    defparam selected_i0.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut_4_lut_adj_697 (.A(selected[0]), .B(selected[1]), 
         .C(LM32D_SEL_O[2]), .D(n18080), .Z(REF_CLK_c_enable_1597)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C (D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam i1_2_lut_4_lut_4_lut_adj_697.init = 16'h6200;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_698 (.A(selected[0]), .B(selected[1]), 
         .C(LM32D_SEL_O[3]), .D(n18080), .Z(REF_CLK_c_enable_1605)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C (D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(321[22:38])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_698.init = 16'h6200;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_699 (.A(selected[0]), .B(selected[1]), 
         .C(LM32D_SEL_O[1]), .D(n18080), .Z(REF_CLK_c_enable_1589)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C (D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(321[22:38])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_699.init = 16'h6200;
    LUT4 i14884_2_lut_rep_924_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[1]), 
         .Z(n41329)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14884_2_lut_rep_924_3_lut.init = 16'h4040;
    LUT4 i1_3_lut_4_lut_adj_700 (.A(selected[0]), .B(selected[1]), .C(locked_N_493), 
         .D(n41387), .Z(n9)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_3_lut_4_lut_adj_700.init = 16'h0040;
    LUT4 i33081_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\counter[2] ), 
         .Z(n12390)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i33081_2_lut_3_lut.init = 16'hbfbf;
    LUT4 i1_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\LM32D_ADR_O[0] ), 
         .Z(n71_adj_305)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h4040;
    LUT4 EBR_DAT_O_15__I_0_i3_3_lut_4_lut (.A(n41429), .B(n41306), .C(\SHAREDBUS_DAT_I[10] ), 
         .D(ebrEBR_DAT_O[10]), .Z(\genblk1.write_data_15__N_3557 [2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam EBR_DAT_O_15__I_0_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_rep_1061 (.A(n45101), .B(selected[0]), .C(\LM32D_ADR_O[6] ), 
         .Z(n45081)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_rep_1061.init = 16'h2020;
    LUT4 i1_3_lut_rep_1056 (.A(selected[1]), .B(selected[0]), .C(\LM32D_ADR_O[12] ), 
         .Z(n45076)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_rep_1056.init = 16'h2020;
    LUT4 WBS_ADR_I_31__I_0_i7_3_lut_rep_941_4_lut_4_lut (.A(selected[1]), 
         .B(selected[0]), .C(\LM32D_ADR_O[6] ), .D(\LM32I_ADR_O[6] ), 
         .Z(n41346)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam WBS_ADR_I_31__I_0_i7_3_lut_rep_941_4_lut_4_lut.init = 16'h6420;
    LUT4 i11097_3_lut_rep_898_4_lut_4_lut (.A(selected[1]), .B(selected[0]), 
         .C(\LM32D_ADR_O[12] ), .D(\LM32I_ADR_O[12] ), .Z(n41303)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam i11097_3_lut_rep_898_4_lut_4_lut.init = 16'h6420;
    LUT4 i1_3_lut_rep_1062 (.A(n45101), .B(n45097), .C(\LM32D_ADR_O[4] ), 
         .Z(n45082)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_rep_1062.init = 16'h2020;
    LUT4 i1_3_lut_rep_1057 (.A(selected[1]), .B(n45097), .C(\LM32D_ADR_O[9] ), 
         .Z(n45077)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_rep_1057.init = 16'h2020;
    LUT4 WBS_ADR_I_31__I_0_i5_3_lut_rep_942_4_lut_4_lut (.A(selected[1]), 
         .B(selected[0]), .C(\LM32D_ADR_O[4] ), .D(\LM32I_ADR_O[4] ), 
         .Z(n41347)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam WBS_ADR_I_31__I_0_i5_3_lut_rep_942_4_lut_4_lut.init = 16'h6420;
    LUT4 WBS_ADR_I_31__I_0_i10_3_lut_rep_905_4_lut_4_lut (.A(selected[1]), 
         .B(selected[0]), .C(\LM32D_ADR_O[9] ), .D(\LM32I_ADR_O[9] ), 
         .Z(n41310)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam WBS_ADR_I_31__I_0_i10_3_lut_rep_905_4_lut_4_lut.init = 16'h6420;
    LUT4 i33065_2_lut_rep_817_4_lut_4_lut_4_lut_4_lut (.A(selected[0]), .B(selected[1]), 
         .C(\LM32D_CTI_O[0] ), .D(\LM32I_CTI_O[0] ), .Z(n41222)) /* synthesis lut_function=(!(A (B+(D))+!A ((C)+!B))) */ ;
    defparam i33065_2_lut_rep_817_4_lut_4_lut_4_lut_4_lut.init = 16'h0426;
    LUT4 i14514_2_lut_rep_899_3_lut (.A(n45097), .B(n45101), .C(LM32D_WE_O), 
         .Z(n41304)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14514_2_lut_rep_899_3_lut.init = 16'h4040;
    LUT4 i2_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(n38693), 
         .Z(n6034)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i2_2_lut_3_lut.init = 16'h4040;
    LUT4 i14885_2_lut_rep_925_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[2]), 
         .Z(n41330)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14885_2_lut_rep_925_3_lut.init = 16'h4040;
    LUT4 i14886_2_lut_rep_926_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[3]), 
         .Z(n41331)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14886_2_lut_rep_926_3_lut.init = 16'h4040;
    LUT4 i14887_2_lut_rep_927_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[4]), 
         .Z(n41332)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14887_2_lut_rep_927_3_lut.init = 16'h4040;
    LUT4 i14888_2_lut_rep_928_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[5]), 
         .Z(n41333)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14888_2_lut_rep_928_3_lut.init = 16'h4040;
    LUT4 i14889_2_lut_rep_929_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[6]), 
         .Z(n41334)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14889_2_lut_rep_929_3_lut.init = 16'h4040;
    LUT4 i14890_2_lut_rep_930_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[7]), 
         .Z(n41335)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14890_2_lut_rep_930_3_lut.init = 16'h4040;
    LUT4 i14899_2_lut_rep_931_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[16]), 
         .Z(n41336)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14899_2_lut_rep_931_3_lut.init = 16'h4040;
    LUT4 i14900_2_lut_rep_932_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[17]), 
         .Z(n41337)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14900_2_lut_rep_932_3_lut.init = 16'h4040;
    LUT4 i14901_2_lut_rep_933_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[18]), 
         .Z(n41338)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14901_2_lut_rep_933_3_lut.init = 16'h4040;
    LUT4 i14902_2_lut_rep_934_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[19]), 
         .Z(n41339)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14902_2_lut_rep_934_3_lut.init = 16'h4040;
    LUT4 EBR_DAT_O_15__I_0_i2_3_lut_4_lut (.A(n41429), .B(n41306), .C(\SHAREDBUS_DAT_I[9] ), 
         .D(ebrEBR_DAT_O[9]), .Z(\genblk1.write_data_15__N_3557 [1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam EBR_DAT_O_15__I_0_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4857_2_lut_3_lut_4_lut (.A(n41429), .B(n41306), .C(n41278), 
         .D(n41193), .Z(REF_CLK_c_enable_1558)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam i4857_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i14903_2_lut_rep_935_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[20]), 
         .Z(n41340)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14903_2_lut_rep_935_3_lut.init = 16'h4040;
    LUT4 i14904_2_lut_rep_936_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[21]), 
         .Z(n41341)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14904_2_lut_rep_936_3_lut.init = 16'h4040;
    LUT4 i14905_2_lut_rep_937_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[22]), 
         .Z(n41342)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14905_2_lut_rep_937_3_lut.init = 16'h4040;
    LUT4 i14906_2_lut_rep_938_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_DAT_O[23]), 
         .Z(n41343)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i14906_2_lut_rep_938_3_lut.init = 16'h4040;
    LUT4 mux_9_i4_3_lut_4_lut (.A(n41429), .B(n41307), .C(\SHAREDBUS_DAT_I[27] ), 
         .D(data[27]), .Z(n96[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_9_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4682_3_lut_4_lut_then_4_lut (.A(\LM32D_ADR_O[7] ), .B(selected[0]), 
         .C(selected[1]), .D(n55), .Z(n41484)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (B (D)+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i4682_3_lut_4_lut_then_4_lut.init = 16'hef20;
    LUT4 mux_9_i1_3_lut_4_lut (.A(n41429), .B(n41307), .C(\SHAREDBUS_DAT_I[24] ), 
         .D(data[24]), .Z(n96[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_9_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4682_3_lut_4_lut_else_4_lut (.A(n55), .Z(n41483)) /* synthesis lut_function=(A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i4682_3_lut_4_lut_else_4_lut.init = 16'haaaa;
    LUT4 mux_9_i5_3_lut_4_lut (.A(n41429), .B(n41307), .C(\SHAREDBUS_DAT_I[28] ), 
         .D(data[28]), .Z(n96[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_9_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 LM32D_SEL_O_1__bdd_4_lut (.A(LM32D_SEL_O[1]), .B(LM32D_SEL_O[3]), 
         .C(LM32D_SEL_O[2]), .D(LM32D_SEL_O[0]), .Z(n38693)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B (C+(D))+!B (C (D)+!C !(D))))) */ ;
    defparam LM32D_SEL_O_1__bdd_4_lut.init = 16'h0116;
    LUT4 mux_9_i6_3_lut_4_lut (.A(n41429), .B(n41307), .C(\SHAREDBUS_DAT_I[29] ), 
         .D(data[29]), .Z(n96[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_9_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_4_lut_adj_701 (.A(n41429), .B(n41307), .C(n41304), .D(n41279), 
         .Z(n29830)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam i1_3_lut_4_lut_adj_701.init = 16'h00e0;
    LUT4 mux_9_i3_3_lut_4_lut (.A(n41429), .B(n41307), .C(\SHAREDBUS_DAT_I[26] ), 
         .D(data[26]), .Z(n96[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_9_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i2_3_lut_4_lut (.A(n41429), .B(n41307), .C(\SHAREDBUS_DAT_I[25] ), 
         .D(data[25]), .Z(n96[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_9_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4889_2_lut_3_lut_4_lut (.A(n41429), .B(n41307), .C(n41278), 
         .D(n41193), .Z(REF_CLK_c_enable_1574)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam i4889_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 EBR_DAT_O_31__I_0_i3_3_lut_4_lut (.A(n41429), .B(n41307), .C(\SHAREDBUS_DAT_I[26] ), 
         .D(ebrEBR_DAT_O[26]), .Z(\genblk1.write_data_31__N_3525 [2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam EBR_DAT_O_31__I_0_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i7_3_lut_4_lut (.A(n41429), .B(n41307), .C(\SHAREDBUS_DAT_I[30] ), 
         .D(data[30]), .Z(n96[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_9_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 EBR_DAT_O_31__I_0_i8_3_lut_4_lut (.A(n41429), .B(n41307), .C(\SHAREDBUS_DAT_I[31] ), 
         .D(ebrEBR_DAT_O[31]), .Z(\genblk1.write_data_31__N_3525 [7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam EBR_DAT_O_31__I_0_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 EBR_DAT_O_31__I_0_i7_3_lut_4_lut (.A(n41429), .B(n41307), .C(\SHAREDBUS_DAT_I[30] ), 
         .D(ebrEBR_DAT_O[30]), .Z(\genblk1.write_data_31__N_3525 [6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam EBR_DAT_O_31__I_0_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 EBR_DAT_O_31__I_0_i6_3_lut_4_lut (.A(n41429), .B(n41307), .C(\SHAREDBUS_DAT_I[29] ), 
         .D(ebrEBR_DAT_O[29]), .Z(\genblk1.write_data_31__N_3525 [5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam EBR_DAT_O_31__I_0_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 EBR_DAT_O_31__I_0_i5_3_lut_4_lut (.A(n41429), .B(n41307), .C(\SHAREDBUS_DAT_I[28] ), 
         .D(ebrEBR_DAT_O[28]), .Z(\genblk1.write_data_31__N_3525 [4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam EBR_DAT_O_31__I_0_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_9_i8_3_lut_4_lut (.A(n41429), .B(n41307), .C(\SHAREDBUS_DAT_I[31] ), 
         .D(data[31]), .Z(n96[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam mux_9_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 EBR_DAT_O_31__I_0_i4_3_lut_4_lut (.A(n41429), .B(n41307), .C(\SHAREDBUS_DAT_I[27] ), 
         .D(ebrEBR_DAT_O[27]), .Z(\genblk1.write_data_31__N_3525 [3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam EBR_DAT_O_31__I_0_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 EBR_DAT_O_31__I_0_i2_3_lut_4_lut (.A(n41429), .B(n41307), .C(\SHAREDBUS_DAT_I[25] ), 
         .D(ebrEBR_DAT_O[25]), .Z(\genblk1.write_data_31__N_3525 [1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam EBR_DAT_O_31__I_0_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 EBR_DAT_O_31__I_0_i1_3_lut_4_lut (.A(n41429), .B(n41307), .C(\SHAREDBUS_DAT_I[24] ), 
         .D(ebrEBR_DAT_O[24]), .Z(\genblk1.write_data_31__N_3525 [0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam EBR_DAT_O_31__I_0_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_9_i3_2_lut_rep_981 (.A(selected[0]), .B(selected[1]), .Z(n41386)) /* synthesis lut_function=(A+(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(253[7:20])
    defparam equal_9_i3_2_lut_rep_981.init = 16'heeee;
    LUT4 i1_3_lut_rep_900_4_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_STB_O), 
         .D(\selected_1__N_354[0] ), .Z(REF_CLK_c_enable_1623)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(253[7:20])
    defparam i1_3_lut_rep_900_4_lut.init = 16'hfffe;
    PFUMX i34373 (.BLUT(n41480), .ALUT(n41481), .C0(LM32D_WE_O), .Z(n41482));
    LUT4 i14512_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\selected_1__N_354[0] ), 
         .Z(selected_1__N_350[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(253[7:20])
    defparam i14512_2_lut_3_lut.init = 16'h1010;
    LUT4 i31169_4_lut_4_lut (.A(selected[0]), .B(selected[1]), .C(n9234), 
         .D(\selected_1__N_354[0] ), .Z(n36341)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(253[7:20])
    defparam i31169_4_lut_4_lut.init = 16'h0c1d;
    LUT4 selected_1__I_0_91_i3_2_lut_rep_985 (.A(selected[0]), .B(selected[1]), 
         .Z(n41390)) /* synthesis lut_function=((B)+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam selected_1__I_0_91_i3_2_lut_rep_985.init = 16'hdddd;
    LUT4 i1_3_lut_4_lut_adj_702 (.A(selected[0]), .B(selected[1]), .C(\next_cycle_type[2] ), 
         .D(\LM32I_ADR_O[2] ), .Z(n32216)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam i1_3_lut_4_lut_adj_702.init = 16'hdfff;
    LUT4 i4678_3_lut_4_lut_then_4_lut (.A(\LM32D_ADR_O[5] ), .B(selected[0]), 
         .C(selected[1]), .D(n61_adj_306), .Z(n41487)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (B (D)+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i4678_3_lut_4_lut_then_4_lut.init = 16'hef20;
    LUT4 i4678_3_lut_4_lut_else_4_lut (.A(n61_adj_306), .Z(n41486)) /* synthesis lut_function=(A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i4678_3_lut_4_lut_else_4_lut.init = 16'haaaa;
    LUT4 i14795_3_lut_rep_851_4_lut (.A(selected[0]), .B(selected[1]), .C(n21), 
         .D(n33), .Z(n41256)) /* synthesis lut_function=(A (B ((D)+!C))+!A ((D)+!C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(316[22:38])
    defparam i14795_3_lut_rep_851_4_lut.init = 16'hdd0d;
    LUT4 i1_2_lut (.A(n31955), .B(n953[0]), .Z(n32220)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut.init = 16'h4444;
    FD1P3DX selected_i1_rep_1067 (.D(n36341), .SP(REF_CLK_c_enable_1623), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(n45101)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=1, LSE_RCOL=20, LSE_LLINE=488, LSE_RLINE=529 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(252[7] 275[5])
    defparam selected_i1_rep_1067.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n34850), .B(n41210), .C(n15_adj_307), .D(n35868), 
         .Z(n18080)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i1_4_lut.init = 16'h0008;
    LUT4 i1_4_lut_adj_703 (.A(n34836), .B(n41225), .C(n19), .D(n41226), 
         .Z(n34850)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i1_4_lut_adj_703.init = 16'h0200;
    LUT4 i1_4_lut_adj_704 (.A(\SHAREDBUS_ADR_I[30] ), .B(n41260), .C(n41278), 
         .D(n34816), .Z(n34836)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i1_4_lut_adj_704.init = 16'h1000;
    LUT4 i1_3_lut_4_lut_3_lut_4_lut (.A(n45097), .B(n45101), .C(LM32D_SEL_O[0]), 
         .D(LM32D_SEL_O[1]), .Z(n11831)) /* synthesis lut_function=(A (B)+!A !(B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(321[22:38])
    defparam i1_3_lut_4_lut_3_lut_4_lut.init = 16'h9ddd;
    LUT4 selected_1__I_0_i3_2_lut_rep_1022 (.A(selected[0]), .B(selected[1]), 
         .Z(n41427)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(321[22:38])
    defparam selected_1__I_0_i3_2_lut_rep_1022.init = 16'hbbbb;
    LUT4 i15508_2_lut_rep_918_3_lut_2_lut (.A(selected[0]), .B(n45101), 
         .Z(n41323)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(321[22:38])
    defparam i15508_2_lut_rep_918_3_lut_2_lut.init = 16'h9999;
    LUT4 i1_3_lut_4_lut_adj_705 (.A(n45097), .B(n45101), .C(LM32D_SEL_O[3]), 
         .D(LM32D_SEL_O[2]), .Z(n33)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(321[22:38])
    defparam i1_3_lut_4_lut_adj_705.init = 16'hbfff;
    LUT4 i1_2_lut_rep_1024 (.A(n45097), .B(n45101), .Z(n41429)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_1024.init = 16'h2222;
    LUT4 i1_3_lut_rep_904_4_lut_3_lut (.A(n45097), .B(n45101), .C(LM32D_SEL_O[2]), 
         .Z(n41309)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;
    defparam i1_3_lut_rep_904_4_lut_3_lut.init = 16'h6262;
    LUT4 i1_2_lut_rep_834_3_lut_4_lut_3_lut (.A(selected[0]), .B(selected[1]), 
         .C(LM32D_SEL_O[3]), .Z(n41239)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;
    defparam i1_2_lut_rep_834_3_lut_4_lut_3_lut.init = 16'h6262;
    LUT4 i1_2_lut_rep_833_3_lut_4_lut_3_lut (.A(selected[0]), .B(selected[1]), 
         .C(LM32D_SEL_O[1]), .Z(n41238)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;
    defparam i1_2_lut_rep_833_3_lut_4_lut_3_lut.init = 16'h6262;
    LUT4 i1_2_lut_rep_765_3_lut_4_lut (.A(selected[0]), .B(selected[1]), 
         .C(n13990), .D(bus_error_f_N_1884), .Z(REF_CLK_c_enable_1131)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_rep_765_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_3_lut_rep_919_4_lut_3_lut (.A(n45097), .B(n45101), .C(LM32D_SEL_O[0]), 
         .Z(n41324)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;
    defparam i1_3_lut_rep_919_4_lut_3_lut.init = 16'h6262;
    LUT4 i1_2_lut_rep_816_4_lut_4_lut_4_lut_4_lut (.A(selected[0]), .B(selected[1]), 
         .C(\LM32D_CTI_O[0] ), .D(\LM32I_CTI_O[0] ), .Z(n41221)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)))) */ ;
    defparam i1_2_lut_rep_816_4_lut_4_lut_4_lut_4_lut.init = 16'h6240;
    LUT4 i1_3_lut_rep_1051 (.A(n45101), .B(n45097), .C(\LM32D_ADR_O[14] ), 
         .Z(n45071)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_rep_1051.init = 16'h2020;
    LUT4 WBS_ADR_I_31__I_0_i15_3_lut_rep_893_4_lut_4_lut (.A(selected[1]), 
         .B(selected[0]), .C(\LM32D_ADR_O[14] ), .D(\LM32I_ADR_O[14] ), 
         .Z(n41298)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam WBS_ADR_I_31__I_0_i15_3_lut_rep_893_4_lut_4_lut.init = 16'h6420;
    LUT4 i4224_2_lut_3_lut_4_lut (.A(n41304), .B(write_ack), .C(n41324), 
         .D(n41193), .Z(REF_CLK_c_enable_1550)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i4224_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i4873_2_lut_3_lut_4_lut (.A(n41304), .B(write_ack), .C(n41309), 
         .D(n41193), .Z(REF_CLK_c_enable_1566)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(292[2] 293[4])
    defparam i4873_2_lut_3_lut_4_lut.init = 16'h2000;
    PFUMX i35861 (.BLUT(n45083), .ALUT(n45084), .C0(\LM32I_CTI_O[0] ), 
          .Z(n9234));
    LUT4 i1_3_lut_rep_1059 (.A(n45101), .B(n45097), .C(\LM32D_ADR_O[2] ), 
         .Z(n45079)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_rep_1059.init = 16'h2020;
    LUT4 i1_3_lut_rep_1052 (.A(selected[1]), .B(selected[0]), .C(\LM32D_ADR_O[13] ), 
         .Z(n45072)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_rep_1052.init = 16'h2020;
    LUT4 i8684_3_lut_rep_940_4_lut_4_lut (.A(n45101), .B(n45097), .C(\LM32D_ADR_O[2] ), 
         .D(\LM32I_ADR_O[2] ), .Z(n41345)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam i8684_3_lut_rep_940_4_lut_4_lut.init = 16'h6420;
    LUT4 WBS_ADR_I_31__I_0_i14_3_lut_rep_895_4_lut_4_lut (.A(n45101), .B(n45097), 
         .C(\LM32D_ADR_O[13] ), .D(\LM32I_ADR_O[13] ), .Z(n41300)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam WBS_ADR_I_31__I_0_i14_3_lut_rep_895_4_lut_4_lut.init = 16'h6420;
    LUT4 i1_3_lut_rep_1060 (.A(n45101), .B(n45097), .C(\next_cycle_type[2]_adj_308 ), 
         .Z(n45080)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_rep_1060.init = 16'h2020;
    LUT4 i1_3_lut_rep_1053 (.A(selected[1]), .B(selected[0]), .C(\LM32D_ADR_O[11] ), 
         .Z(n45073)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_rep_1053.init = 16'h2020;
    LUT4 i8683_rep_141_3_lut_4_lut_4_lut (.A(selected[1]), .B(selected[0]), 
         .C(\next_cycle_type[2]_adj_308 ), .D(\next_cycle_type[2] ), .Z(n37905)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam i8683_rep_141_3_lut_4_lut_4_lut.init = 16'h6420;
    LUT4 WBS_ADR_I_31__I_0_i12_3_lut_rep_894_4_lut_4_lut (.A(selected[1]), 
         .B(n45097), .C(\LM32D_ADR_O[11] ), .D(\LM32I_ADR_O[11] ), .Z(n41299)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam WBS_ADR_I_31__I_0_i12_3_lut_rep_894_4_lut_4_lut.init = 16'h6420;
    LUT4 i8683_rep_140_3_lut_4_lut_4_lut (.A(selected[1]), .B(selected[0]), 
         .C(\next_cycle_type[2]_adj_308 ), .D(\next_cycle_type[2] ), .Z(n37904)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam i8683_rep_140_3_lut_4_lut_4_lut.init = 16'h6420;
    LUT4 i1_3_lut_rep_1054 (.A(n45101), .B(n45097), .C(\LM32D_ADR_O[8] ), 
         .Z(n45074)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_rep_1054.init = 16'h2020;
    LUT4 i8683_rep_142_3_lut_4_lut_4_lut (.A(selected[1]), .B(selected[0]), 
         .C(\next_cycle_type[2]_adj_308 ), .D(\next_cycle_type[2] ), .Z(n37906)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam i8683_rep_142_3_lut_4_lut_4_lut.init = 16'h6420;
    LUT4 WBS_ADR_I_31__I_0_i9_3_lut_rep_896_4_lut_4_lut (.A(selected[1]), 
         .B(selected[0]), .C(\LM32D_ADR_O[8] ), .D(\LM32I_ADR_O[8] ), 
         .Z(n41301)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam WBS_ADR_I_31__I_0_i9_3_lut_rep_896_4_lut_4_lut.init = 16'h6420;
    LUT4 i8683_3_lut_rep_939_4_lut_4_lut (.A(selected[1]), .B(selected[0]), 
         .C(\next_cycle_type[2]_adj_308 ), .D(\next_cycle_type[2] ), .Z(n41344)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam i8683_3_lut_rep_939_4_lut_4_lut.init = 16'h6420;
    LUT4 i8683_rep_139_3_lut_4_lut_4_lut (.A(selected[1]), .B(selected[0]), 
         .C(\next_cycle_type[2]_adj_308 ), .D(\next_cycle_type[2] ), .Z(n37903)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;
    defparam i8683_rep_139_3_lut_4_lut_4_lut.init = 16'h6420;
    
endmodule
//
// Verilog Description of module lm32_top
//

module lm32_top (GND_net, n41300, n41194, LEDGPIO_ACK_O, n1128, REF_CLK_c, 
            n69, REF_CLK_c_enable_1606, \state_1__N_3407[1] , ROM_DAT_O, 
            write_enable, n6362, n78, n87, n96, \counter[2] , n41246, 
            n19808, data, \SHAREDBUS_ADR_I[10] , n41310, n41301, \SHAREDBUS_ADR_I[7] , 
            n41346, \SHAREDBUS_ADR_I[5] , n41347, n41344, n41345, 
            VCC_net, write_idx_w, n41352, n41351, w_result, n41350, 
            dcache_refill_request, \operand_1_x[1] , dc_re, n41430, 
            n41432, REF_CLK_c_enable_176, n7611, n41405, REF_CLK_c_enable_164, 
            n41380, LM32D_CYC_O, locked_N_493, n41356, n41355, n41353, 
            n41358, n41359, \operand_m[10] , \operand_m[9] , \operand_m[5] , 
            LM32D_WE_O, dcache_select_x, n31750, n31955, n30241, n953, 
            n41326, n41354, bie, n31279, \adder_result_x[16] , \adder_result_x[17] , 
            \adder_result_x[18] , \adder_result_x[19] , \adder_result_x[20] , 
            \adder_result_x[21] , \adder_result_x[22] , \adder_result_x[23] , 
            \adder_result_x[24] , \adder_result_x[25] , \adder_result_x[26] , 
            \adder_result_x[27] , \adder_result_x[28] , \adder_result_x[29] , 
            \adder_result_x[30] , \adder_result_x[31] , n6518, n6648, 
            bus_error_f_N_1884, branch_target_d, direction_m, n45103, 
            n45099, n41394, n41401, bie_N_3274, pc_f, n41325, n17816, 
            n41379, \shifter_result_m[21] , n41357, \left_shift_result[21] , 
            \left_shift_result[10] , b, \p[0] , \p[1] , \p[2] , \p[3] , 
            \p[4] , \p[5] , \p[6] , \p[7] , \p[8] , \p[9] , \p[10] , 
            \p[11] , \p[12] , \p[13] , \p[14] , \p[15] , \p[16] , 
            \p[17] , \p[18] , \p[19] , \p[20] , \p[21] , \p[22] , 
            \p[23] , \p[24] , \p[25] , \p[26] , \p[27] , \p[28] , 
            \p[29] , \p[30] , \a[31] , t, LM32D_DAT_O, REF_CLK_c_enable_1221, 
            SHAREDBUS_DAT_O, LM32D_SEL_O, \LM32D_ADR_O[0] , \LM32D_CTI_O[0] , 
            n38965, LM32D_STB_O, n21, \LM32D_ADR_O[1] , \LM32D_ADR_O[2] , 
            \next_cycle_type[2] , \LM32D_ADR_O[4] , \LM32D_ADR_O[5] , 
            \d_adr_o_31__N_2278[5] , \LM32D_ADR_O[6] , \LM32D_ADR_O[7] , 
            \LM32D_ADR_O[8] , \LM32D_ADR_O[9] , \d_adr_o_31__N_2278[9] , 
            \LM32D_ADR_O[10] , \d_adr_o_31__N_2278[10] , \LM32D_ADR_O[11] , 
            \LM32D_ADR_O[12] , \LM32D_ADR_O[13] , \LM32D_ADR_O[14] , \LM32D_ADR_O[15] , 
            \LM32D_ADR_O[16] , \LM32D_ADR_O[17] , \LM32D_ADR_O[18] , \LM32D_ADR_O[19] , 
            \LM32D_ADR_O[20] , \LM32D_ADR_O[21] , \LM32D_ADR_O[22] , \LM32D_ADR_O[23] , 
            \LM32D_ADR_O[24] , \LM32D_ADR_O[25] , \LM32D_ADR_O[26] , \LM32D_ADR_O[27] , 
            \LM32D_ADR_O[28] , \LM32D_ADR_O[29] , \LM32D_ADR_O[30] , \LM32D_ADR_O[31] , 
            n41387, n9, \state[0] , \state[2] , flush_set, flush_set_8__N_2513, 
            \dcache_refill_address[5] , \dcache_refill_address[9] , \dcache_refill_address[10] , 
            \tmem_write_address[1] , \tmem_write_address[5] , \tmem_write_address[6] , 
            \dmem_write_address[3] , \dmem_write_address[7] , \dmem_write_address[8] , 
            n36337, SPI_INT_O_N_4422, SPI_INT_O_N_4417, SPI_INT_O_N_4421, 
            \genblk1.wait_one_tick_done , n6781, n6764, n6749, n41410, 
            n13990, n32216, \LM32I_CTI_O[0] , REF_CLK_c_enable_97, n30900, 
            pc_d, REF_CLK_c_enable_1131, n6760, n45105, n73_adj_232, 
            n41461, \next_cycle_type[2]_adj_233 , n45080, n41390, n5223, 
            n37955, n37956, n37954, n41250, n41251, n41279, \LM32I_ADR_O[2] , 
            n45079, \reg_12[2] , n2, \reg_12[12] , n40677, \reg_12[29] , 
            n2_adj_234, \reg_12[3] , n2_adj_235, \reg_12[6] , n2_adj_236, 
            \reg_12[4] , n2_adj_237, \reg_12[14] , n2_adj_238, n41429, 
            \reg_12[22] , n2_adj_239, \reg_12[13] , n2_adj_240, \reg_12[21] , 
            n2_adj_241, \reg_12[28] , n2_adj_242, \reg_12[11] , n2_adj_243, 
            \reg_12[18] , n2_adj_244, \reg_12[25] , n2_adj_245, \reg_12[9] , 
            n2_adj_246, \reg_12[17] , n2_adj_247, \reg_12[24] , n2_adj_248, 
            \reg_12[7] , n2_adj_249, \reg_12[15] , n2_adj_250, n6589, 
            n6584, n37179, n6439, n6434, n37177, n6599, n6594, 
            n37180, n6629, n6624, n37183, n6579, n6574, n37178, 
            n6429, n6424, n37176, n6609, n6604, n37181, n6619, 
            n6614, n37182, n37185, n37184, n37188, n37187, n37186, 
            n37189, n7603, n7571, n7607, n7575, n7606, n7574, 
            n7604, n7572, n7605, n7573, n7608, n7576, n7602, n7570, 
            \selected_1__N_354[0] , n7601, n7569, n7600, n7568, n7599, 
            n7567, n7598, n7566, n7597, n7565, n7596, n7564, n7595, 
            n7563, n7594, n7562, n7593, n7561, n7592, n7560, n7584, 
            n7552, n7583, n7551, n7582, n7550, n7581, n7549, n7580, 
            n7548, n7579, n7547, n7578, n7546, n7577, n7545, n6750, 
            n7591, n7559, n7590, n7558, n7589, n7557, n7588, n7556, 
            n7587, n7555, n7586, n7554, n7585, n7553, n37501, 
            n37500, n37502, n37499, n37498, n37497, n37496, n6751, 
            n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, 
            n6761, n6762, n6763, n37495, n7672, n7640, n7673, 
            n7641, n34, n7674, n7642, n7675, n7643, n7676, n7644, 
            n7671, n7639, n7670, n7638, n7669, n7637, n7668, n7636, 
            n7667, n7635, n7666, n7634, n7665, n7633, n7664, n7632, 
            n7663, n7631, n7662, n7630, n7661, n7629, n7660, n7628, 
            n36, n7652, n7620, n7651, n7619, n7650, n7618, n7649, 
            n7617, n37, n7648, n7616, n7647, n7615, n7646, n7614, 
            n7645, n7613, n7659, n7627, n7658, n7626, n7657, n7625, 
            n7656, n7624, n7655, n7623, n7654, n7622, n7653, n7621, 
            n37504, n37503, n37507, n37506, n37505, n37508, n45106, 
            \LM32I_ADR_O[4] , \LM32I_ADR_O[5] , \LM32I_ADR_O[6] , \LM32I_ADR_O[7] , 
            \LM32I_ADR_O[8] , \LM32I_ADR_O[9] , \LM32I_ADR_O[10] , \LM32I_ADR_O[11] , 
            \LM32I_ADR_O[12] , \LM32I_ADR_O[13] , \LM32I_ADR_O[14] , \LM32I_ADR_O[15] , 
            \LM32I_ADR_O[16] , \LM32I_ADR_O[17] , \LM32I_ADR_O[18] , \LM32I_ADR_O[19] , 
            \LM32I_ADR_O[20] , \LM32I_ADR_O[21] , \LM32I_ADR_O[22] , \LM32I_ADR_O[23] , 
            \LM32I_ADR_O[24] , \LM32I_ADR_O[25] , \LM32I_ADR_O[26] , \LM32I_ADR_O[27] , 
            \LM32I_ADR_O[28] , \LM32I_ADR_O[29] , \LM32I_ADR_O[30] , \LM32I_ADR_O[31] , 
            n949, n32220, selected, flush_set_adj_272, flush_set_8__N_1953, 
            n157, n36336, n10589, n10585, n10591, n10593, n10587, 
            n10595, n10452) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input n41300;
    input n41194;
    input LEDGPIO_ACK_O;
    output n1128;
    input REF_CLK_c;
    input [7:0]n69;
    input REF_CLK_c_enable_1606;
    output \state_1__N_3407[1] ;
    output [31:0]ROM_DAT_O;
    output write_enable;
    input n6362;
    input [7:0]n78;
    input [7:0]n87;
    input [7:0]n96;
    input \counter[2] ;
    input n41246;
    input n19808;
    output [31:0]data;
    input \SHAREDBUS_ADR_I[10] ;
    input n41310;
    input n41301;
    input \SHAREDBUS_ADR_I[7] ;
    input n41346;
    input \SHAREDBUS_ADR_I[5] ;
    input n41347;
    input n41344;
    input n41345;
    input VCC_net;
    output [4:0]write_idx_w;
    output n41352;
    output n41351;
    output [31:0]w_result;
    output n41350;
    output dcache_refill_request;
    output \operand_1_x[1] ;
    output dc_re;
    output n41430;
    input n41432;
    output REF_CLK_c_enable_176;
    output n7611;
    input n41405;
    output REF_CLK_c_enable_164;
    input n41380;
    output LM32D_CYC_O;
    output locked_N_493;
    output n41356;
    output n41355;
    output n41353;
    output n41358;
    output n41359;
    output \operand_m[10] ;
    output \operand_m[9] ;
    output \operand_m[5] ;
    output LM32D_WE_O;
    input dcache_select_x;
    input n31750;
    input n31955;
    input n30241;
    input [0:0]n953;
    input n41326;
    output n41354;
    output bie;
    output n31279;
    output \adder_result_x[16] ;
    output \adder_result_x[17] ;
    output \adder_result_x[18] ;
    output \adder_result_x[19] ;
    output \adder_result_x[20] ;
    output \adder_result_x[21] ;
    output \adder_result_x[22] ;
    output \adder_result_x[23] ;
    output \adder_result_x[24] ;
    output \adder_result_x[25] ;
    output \adder_result_x[26] ;
    output \adder_result_x[27] ;
    output \adder_result_x[28] ;
    output \adder_result_x[29] ;
    output \adder_result_x[30] ;
    output \adder_result_x[31] ;
    input n6518;
    input n6648;
    output bus_error_f_N_1884;
    input [31:2]branch_target_d;
    output direction_m;
    output n45103;
    output n45099;
    output n41394;
    output n41401;
    output bie_N_3274;
    output [31:2]pc_f;
    output n41325;
    input n17816;
    output n41379;
    input \shifter_result_m[21] ;
    output n41357;
    output \left_shift_result[21] ;
    output \left_shift_result[10] ;
    output [31:0]b;
    output \p[0] ;
    output \p[1] ;
    output \p[2] ;
    output \p[3] ;
    output \p[4] ;
    output \p[5] ;
    output \p[6] ;
    output \p[7] ;
    output \p[8] ;
    output \p[9] ;
    output \p[10] ;
    output \p[11] ;
    output \p[12] ;
    output \p[13] ;
    output \p[14] ;
    output \p[15] ;
    output \p[16] ;
    output \p[17] ;
    output \p[18] ;
    output \p[19] ;
    output \p[20] ;
    output \p[21] ;
    output \p[22] ;
    output \p[23] ;
    output \p[24] ;
    output \p[25] ;
    output \p[26] ;
    output \p[27] ;
    output \p[28] ;
    output \p[29] ;
    output \p[30] ;
    output \a[31] ;
    input [32:0]t;
    output [31:0]LM32D_DAT_O;
    input REF_CLK_c_enable_1221;
    input [31:0]SHAREDBUS_DAT_O;
    output [3:0]LM32D_SEL_O;
    output \LM32D_ADR_O[0] ;
    output \LM32D_CTI_O[0] ;
    input n38965;
    output LM32D_STB_O;
    output n21;
    output \LM32D_ADR_O[1] ;
    output \LM32D_ADR_O[2] ;
    output \next_cycle_type[2] ;
    output \LM32D_ADR_O[4] ;
    output \LM32D_ADR_O[5] ;
    input \d_adr_o_31__N_2278[5] ;
    output \LM32D_ADR_O[6] ;
    output \LM32D_ADR_O[7] ;
    output \LM32D_ADR_O[8] ;
    output \LM32D_ADR_O[9] ;
    input \d_adr_o_31__N_2278[9] ;
    output \LM32D_ADR_O[10] ;
    input \d_adr_o_31__N_2278[10] ;
    output \LM32D_ADR_O[11] ;
    output \LM32D_ADR_O[12] ;
    output \LM32D_ADR_O[13] ;
    output \LM32D_ADR_O[14] ;
    output \LM32D_ADR_O[15] ;
    output \LM32D_ADR_O[16] ;
    output \LM32D_ADR_O[17] ;
    output \LM32D_ADR_O[18] ;
    output \LM32D_ADR_O[19] ;
    output \LM32D_ADR_O[20] ;
    output \LM32D_ADR_O[21] ;
    output \LM32D_ADR_O[22] ;
    output \LM32D_ADR_O[23] ;
    output \LM32D_ADR_O[24] ;
    output \LM32D_ADR_O[25] ;
    output \LM32D_ADR_O[26] ;
    output \LM32D_ADR_O[27] ;
    output \LM32D_ADR_O[28] ;
    output \LM32D_ADR_O[29] ;
    output \LM32D_ADR_O[30] ;
    output \LM32D_ADR_O[31] ;
    output n41387;
    input n9;
    output \state[0] ;
    output \state[2] ;
    output [8:0]flush_set;
    input [8:0]flush_set_8__N_2513;
    output \dcache_refill_address[5] ;
    output \dcache_refill_address[9] ;
    output \dcache_refill_address[10] ;
    input \tmem_write_address[1] ;
    input \tmem_write_address[5] ;
    input \tmem_write_address[6] ;
    input \dmem_write_address[3] ;
    input \dmem_write_address[7] ;
    input \dmem_write_address[8] ;
    input n36337;
    input SPI_INT_O_N_4422;
    input SPI_INT_O_N_4417;
    input SPI_INT_O_N_4421;
    output \genblk1.wait_one_tick_done ;
    output n6781;
    output n6764;
    output n6749;
    output n41410;
    input n13990;
    input n32216;
    output \LM32I_CTI_O[0] ;
    input REF_CLK_c_enable_97;
    input n30900;
    output [31:2]pc_d;
    input REF_CLK_c_enable_1131;
    output n6760;
    output n45105;
    input n73_adj_232;
    output n41461;
    output \next_cycle_type[2]_adj_233 ;
    input n45080;
    input n41390;
    input n5223;
    output n37955;
    output n37956;
    output n37954;
    output n41250;
    output n41251;
    output n41279;
    output \LM32I_ADR_O[2] ;
    input n45079;
    input \reg_12[2] ;
    output n2;
    input \reg_12[12] ;
    output n40677;
    input \reg_12[29] ;
    output n2_adj_234;
    input \reg_12[3] ;
    output n2_adj_235;
    input \reg_12[6] ;
    output n2_adj_236;
    input \reg_12[4] ;
    output n2_adj_237;
    input \reg_12[14] ;
    output n2_adj_238;
    input n41429;
    input \reg_12[22] ;
    output n2_adj_239;
    input \reg_12[13] ;
    output n2_adj_240;
    input \reg_12[21] ;
    output n2_adj_241;
    input \reg_12[28] ;
    output n2_adj_242;
    input \reg_12[11] ;
    output n2_adj_243;
    input \reg_12[18] ;
    output n2_adj_244;
    input \reg_12[25] ;
    output n2_adj_245;
    input \reg_12[9] ;
    output n2_adj_246;
    input \reg_12[17] ;
    output n2_adj_247;
    input \reg_12[24] ;
    output n2_adj_248;
    input \reg_12[7] ;
    output n2_adj_249;
    input \reg_12[15] ;
    output n2_adj_250;
    input n6589;
    input n6584;
    output n37179;
    input n6439;
    input n6434;
    output n37177;
    input n6599;
    input n6594;
    output n37180;
    input n6629;
    input n6624;
    output n37183;
    input n6579;
    input n6574;
    output n37178;
    input n6429;
    input n6424;
    output n37176;
    input n6609;
    input n6604;
    output n37181;
    input n6619;
    input n6614;
    output n37182;
    input n37185;
    input n37184;
    output n37188;
    input n37187;
    input n37186;
    output n37189;
    input n7603;
    input n7571;
    input n7607;
    input n7575;
    input n7606;
    input n7574;
    input n7604;
    input n7572;
    input n7605;
    input n7573;
    input n7608;
    input n7576;
    input n7602;
    input n7570;
    output \selected_1__N_354[0] ;
    input n7601;
    input n7569;
    input n7600;
    input n7568;
    input n7599;
    input n7567;
    input n7598;
    input n7566;
    input n7597;
    input n7565;
    input n7596;
    input n7564;
    input n7595;
    input n7563;
    input n7594;
    input n7562;
    input n7593;
    input n7561;
    input n7592;
    input n7560;
    input n7584;
    input n7552;
    input n7583;
    input n7551;
    input n7582;
    input n7550;
    input n7581;
    input n7549;
    input n7580;
    input n7548;
    input n7579;
    input n7547;
    input n7578;
    input n7546;
    input n7577;
    input n7545;
    output n6750;
    input n7591;
    input n7559;
    input n7590;
    input n7558;
    input n7589;
    input n7557;
    input n7588;
    input n7556;
    input n7587;
    input n7555;
    input n7586;
    input n7554;
    input n7585;
    input n7553;
    output n37501;
    output n37500;
    output n37502;
    output n37499;
    output n37498;
    output n37497;
    output n37496;
    output n6751;
    output n6752;
    output n6753;
    output n6754;
    output n6755;
    output n6756;
    output n6757;
    output n6758;
    output n6759;
    output n6761;
    output n6762;
    output n6763;
    output n37495;
    input n7672;
    input n7640;
    input n7673;
    input n7641;
    output n34;
    input n7674;
    input n7642;
    input n7675;
    input n7643;
    input n7676;
    input n7644;
    input n7671;
    input n7639;
    input n7670;
    input n7638;
    input n7669;
    input n7637;
    input n7668;
    input n7636;
    input n7667;
    input n7635;
    input n7666;
    input n7634;
    input n7665;
    input n7633;
    input n7664;
    input n7632;
    input n7663;
    input n7631;
    input n7662;
    input n7630;
    input n7661;
    input n7629;
    input n7660;
    input n7628;
    output n36;
    input n7652;
    input n7620;
    input n7651;
    input n7619;
    input n7650;
    input n7618;
    input n7649;
    input n7617;
    output n37;
    input n7648;
    input n7616;
    input n7647;
    input n7615;
    input n7646;
    input n7614;
    input n7645;
    input n7613;
    input n7659;
    input n7627;
    input n7658;
    input n7626;
    input n7657;
    input n7625;
    input n7656;
    input n7624;
    input n7655;
    input n7623;
    input n7654;
    input n7622;
    input n7653;
    input n7621;
    input n37504;
    input n37503;
    output n37507;
    input n37506;
    input n37505;
    output n37508;
    output n45106;
    output \LM32I_ADR_O[4] ;
    output \LM32I_ADR_O[5] ;
    output \LM32I_ADR_O[6] ;
    output \LM32I_ADR_O[7] ;
    output \LM32I_ADR_O[8] ;
    output \LM32I_ADR_O[9] ;
    output \LM32I_ADR_O[10] ;
    output \LM32I_ADR_O[11] ;
    output \LM32I_ADR_O[12] ;
    output \LM32I_ADR_O[13] ;
    output \LM32I_ADR_O[14] ;
    output \LM32I_ADR_O[15] ;
    output \LM32I_ADR_O[16] ;
    output \LM32I_ADR_O[17] ;
    output \LM32I_ADR_O[18] ;
    output \LM32I_ADR_O[19] ;
    output \LM32I_ADR_O[20] ;
    output \LM32I_ADR_O[21] ;
    output \LM32I_ADR_O[22] ;
    output \LM32I_ADR_O[23] ;
    output \LM32I_ADR_O[24] ;
    output \LM32I_ADR_O[25] ;
    output \LM32I_ADR_O[26] ;
    output \LM32I_ADR_O[27] ;
    output \LM32I_ADR_O[28] ;
    output \LM32I_ADR_O[29] ;
    output \LM32I_ADR_O[30] ;
    output \LM32I_ADR_O[31] ;
    input [0:0]n949;
    input n32220;
    input [1:0]selected;
    output [8:0]flush_set_adj_272;
    input [8:0]flush_set_8__N_1953;
    input [29:0]n157;
    input n36336;
    output n10589;
    output n10585;
    output n10591;
    output n10593;
    output n10587;
    output n10595;
    output n10452;
    
    wire jtag_update /* synthesis is_clock=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(254[6:17])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    wire jtag_update_N_3371 /* synthesis is_inv_clock=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(203[14:23])
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    wire [2:0]jtag_reg_addr_q;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(256[12:27])
    
    wire n41397, jrx_csr_read_data_8__N_3304;
    wire [7:0]jtag_reg_d;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(248[23:33])
    wire [7:0]jtag_reg_q;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(252[12:22])
    wire [2:0]jtag_reg_addr_d;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(255[12:27])
    
    wire rx_toggle_r_r_r, rx_toggle_r_r, n41398, REF_CLK_c_enable_1373, 
        n30162, n41311;
    wire [7:0]uart_tx_byte;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(212[28:40])
    wire [7:0]n4626;
    
    wire n43, n29834, ROM_ACK_O;
    
    LUT4 i1_2_lut_4_lut (.A(jtag_reg_addr_q[2]), .B(n41397), .C(jtag_reg_addr_q[1]), 
         .D(jtag_reg_addr_q[0]), .Z(jrx_csr_read_data_8__N_3304)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0400;
    jtag_cores jtag_cores (.reg_d({jtag_reg_d}), .reg_addr_d({GND_net, jtag_reg_addr_d[1:0]}), 
            .reg_update(jtag_update), .reg_q({jtag_reg_q}), .reg_addr_q({jtag_reg_addr_q})) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=572, LSE_RLINE=613 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(418[12] 432[6])
    LUT4 i15_2_lut_rep_992 (.A(rx_toggle_r_r_r), .B(rx_toggle_r_r), .Z(n41397)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(205[14:27])
    defparam i15_2_lut_rep_992.init = 16'h6666;
    LUT4 i1_2_lut_3_lut (.A(rx_toggle_r_r_r), .B(rx_toggle_r_r), .C(n41398), 
         .Z(REF_CLK_c_enable_1373)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(205[14:27])
    defparam i1_2_lut_3_lut.init = 16'h6060;
    LUT4 i1_3_lut_4_lut (.A(rx_toggle_r_r_r), .B(rx_toggle_r_r), .C(jtag_reg_addr_q[0]), 
         .D(jtag_reg_addr_q[2]), .Z(n30162)) /* synthesis lut_function=(A (B+(C+(D)))+!A ((C+(D))+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(205[14:27])
    defparam i1_3_lut_4_lut.init = 16'hfff9;
    LUT4 i1_3_lut_rep_906_4_lut (.A(rx_toggle_r_r_r), .B(rx_toggle_r_r), 
         .C(jtag_reg_addr_q[1]), .D(jtag_reg_addr_q[2]), .Z(n41311)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A ((C+(D))+!B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(205[14:27])
    defparam i1_3_lut_rep_906_4_lut.init = 16'h0006;
    LUT4 i2_3_lut_rep_993 (.A(jtag_reg_addr_q[0]), .B(jtag_reg_addr_q[2]), 
         .C(jtag_reg_addr_q[1]), .Z(n41398)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(418[12] 432[6])
    defparam i2_3_lut_rep_993.init = 16'h1010;
    LUT4 i1_2_lut_4_lut_adj_646 (.A(jtag_reg_addr_q[0]), .B(jtag_reg_addr_q[2]), 
         .C(jtag_reg_addr_q[1]), .D(uart_tx_byte[0]), .Z(n4626[0])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(418[12] 432[6])
    defparam i1_2_lut_4_lut_adj_646.init = 16'h1000;
    LUT4 i1_2_lut_4_lut_adj_647 (.A(jtag_reg_addr_q[0]), .B(jtag_reg_addr_q[2]), 
         .C(jtag_reg_addr_q[1]), .D(uart_tx_byte[1]), .Z(n4626[1])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(418[12] 432[6])
    defparam i1_2_lut_4_lut_adj_647.init = 16'h1000;
    LUT4 i1_2_lut_4_lut_adj_648 (.A(jtag_reg_addr_q[0]), .B(jtag_reg_addr_q[2]), 
         .C(jtag_reg_addr_q[1]), .D(uart_tx_byte[2]), .Z(n4626[2])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(418[12] 432[6])
    defparam i1_2_lut_4_lut_adj_648.init = 16'h1000;
    LUT4 i1_2_lut_4_lut_adj_649 (.A(jtag_reg_addr_q[0]), .B(jtag_reg_addr_q[2]), 
         .C(jtag_reg_addr_q[1]), .D(uart_tx_byte[3]), .Z(n4626[3])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(418[12] 432[6])
    defparam i1_2_lut_4_lut_adj_649.init = 16'h1000;
    LUT4 i1_2_lut_4_lut_adj_650 (.A(jtag_reg_addr_q[0]), .B(jtag_reg_addr_q[2]), 
         .C(jtag_reg_addr_q[1]), .D(uart_tx_byte[4]), .Z(n4626[4])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(418[12] 432[6])
    defparam i1_2_lut_4_lut_adj_650.init = 16'h1000;
    LUT4 i1_2_lut_4_lut_adj_651 (.A(jtag_reg_addr_q[0]), .B(jtag_reg_addr_q[2]), 
         .C(jtag_reg_addr_q[1]), .D(uart_tx_byte[5]), .Z(n4626[5])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(418[12] 432[6])
    defparam i1_2_lut_4_lut_adj_651.init = 16'h1000;
    LUT4 i1_2_lut_4_lut_adj_652 (.A(jtag_reg_addr_q[0]), .B(jtag_reg_addr_q[2]), 
         .C(jtag_reg_addr_q[1]), .D(uart_tx_byte[6]), .Z(n4626[6])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(418[12] 432[6])
    defparam i1_2_lut_4_lut_adj_652.init = 16'h1000;
    LUT4 i1_2_lut_4_lut_adj_653 (.A(jtag_reg_addr_q[0]), .B(jtag_reg_addr_q[2]), 
         .C(jtag_reg_addr_q[1]), .D(uart_tx_byte[7]), .Z(n4626[7])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(418[12] 432[6])
    defparam i1_2_lut_4_lut_adj_653.init = 16'h1000;
    LUT4 i1_2_lut (.A(jtag_reg_q[5]), .B(jtag_reg_q[6]), .Z(n43)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(418[12] 432[6])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_4_lut (.A(n41311), .B(jtag_reg_addr_q[0]), .C(n43), .D(jtag_reg_q[7]), 
         .Z(n29834)) /* synthesis lut_function=(A (B+!((D)+!C))) */ ;
    defparam i1_4_lut.init = 16'h88a8;
    LUT4 mux_64_i1_4_lut_4_lut (.A(n41300), .B(n41194), .C(ROM_ACK_O), 
         .D(LEDGPIO_ACK_O), .Z(n1128)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(539[44] 547[3])
    defparam mux_64_i1_4_lut_4_lut.init = 16'hdc10;
    INV i35875 (.A(jtag_update), .Z(jtag_update_N_3371));
    lm32_monitor debug_rom (.REF_CLK_c(REF_CLK_c), .n69({n69}), .ROM_ACK_O(ROM_ACK_O), 
            .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), .state_1__N_3407({\state_1__N_3407[1] , 
            Open_8}), .ROM_DAT_O({ROM_DAT_O}), .write_enable(write_enable), 
            .n6362(n6362), .n78({n78}), .n87({n87}), .n96({n96}), .\counter[2] (\counter[2] ), 
            .n41246(n41246), .n19808(n19808), .data({data}), .GND_net(GND_net), 
            .\SHAREDBUS_ADR_I[10] (\SHAREDBUS_ADR_I[10] ), .n41310(n41310), 
            .n41301(n41301), .\SHAREDBUS_ADR_I[7] (\SHAREDBUS_ADR_I[7] ), 
            .n41346(n41346), .\SHAREDBUS_ADR_I[5] (\SHAREDBUS_ADR_I[5] ), 
            .n41347(n41347), .n41344(n41344), .n41345(n41345), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(398[17] 413[8])
    lm32_cpu cpu (.write_idx_w({write_idx_w}), .n41352(n41352), .n41351(n41351), 
            .w_result({w_result}), .n41350(n41350), .REF_CLK_c(REF_CLK_c), 
            .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), .dcache_refill_request(dcache_refill_request), 
            .\operand_1_x[1] (\operand_1_x[1] ), .dc_re(dc_re), .n41430(n41430), 
            .\counter[2] (\counter[2] ), .n41432(n41432), .REF_CLK_c_enable_176(REF_CLK_c_enable_176), 
            .GND_net(GND_net), .n7611(n7611), .n41405(n41405), .REF_CLK_c_enable_164(REF_CLK_c_enable_164), 
            .n41380(n41380), .LM32D_CYC_O(LM32D_CYC_O), .locked_N_493(locked_N_493), 
            .n41356(n41356), .n41355(n41355), .n41353(n41353), .n41358(n41358), 
            .n41359(n41359), .\operand_m[10] (\operand_m[10] ), .\operand_m[9] (\operand_m[9] ), 
            .\operand_m[5] (\operand_m[5] ), .LM32D_WE_O(LM32D_WE_O), .dcache_select_x(dcache_select_x), 
            .n31750(n31750), .n31955(n31955), .n30241(n30241), .n953({n953}), 
            .n41326(n41326), .n41354(n41354), .bie(bie), .n31279(n31279), 
            .\adder_result_x[16] (\adder_result_x[16] ), .\adder_result_x[17] (\adder_result_x[17] ), 
            .\adder_result_x[18] (\adder_result_x[18] ), .\adder_result_x[19] (\adder_result_x[19] ), 
            .\adder_result_x[20] (\adder_result_x[20] ), .\adder_result_x[21] (\adder_result_x[21] ), 
            .\adder_result_x[22] (\adder_result_x[22] ), .\adder_result_x[23] (\adder_result_x[23] ), 
            .\adder_result_x[24] (\adder_result_x[24] ), .\adder_result_x[25] (\adder_result_x[25] ), 
            .\adder_result_x[26] (\adder_result_x[26] ), .\adder_result_x[27] (\adder_result_x[27] ), 
            .\adder_result_x[28] (\adder_result_x[28] ), .\adder_result_x[29] (\adder_result_x[29] ), 
            .\adder_result_x[30] (\adder_result_x[30] ), .\adder_result_x[31] (\adder_result_x[31] ), 
            .n6518(n6518), .n6648(n6648), .bus_error_f_N_1884(bus_error_f_N_1884), 
            .branch_target_d({branch_target_d}), .direction_m(direction_m), 
            .n45103(n45103), .n45099(n45099), .n41394(n41394), .n41401(n41401), 
            .bie_N_3274(bie_N_3274), .pc_f({pc_f}), .VCC_net(VCC_net), 
            .n41325(n41325), .n17816(n17816), .n41379(n41379), .\shifter_result_m[21] (\shifter_result_m[21] ), 
            .\jtag_reg_addr_d[0] (jtag_reg_addr_d[0]), .\jtag_reg_addr_d[1] (jtag_reg_addr_d[1]), 
            .n41357(n41357), .\left_shift_result[21] (\left_shift_result[21] ), 
            .\left_shift_result[10] (\left_shift_result[10] ), .b({b}), 
            .\p[0] (\p[0] ), .\p[1] (\p[1] ), .\p[2] (\p[2] ), .\p[3] (\p[3] ), 
            .\p[4] (\p[4] ), .\p[5] (\p[5] ), .\p[6] (\p[6] ), .\p[7] (\p[7] ), 
            .\p[8] (\p[8] ), .\p[9] (\p[9] ), .\p[10] (\p[10] ), .\p[11] (\p[11] ), 
            .\p[12] (\p[12] ), .\p[13] (\p[13] ), .\p[14] (\p[14] ), .\p[15] (\p[15] ), 
            .\p[16] (\p[16] ), .\p[17] (\p[17] ), .\p[18] (\p[18] ), .\p[19] (\p[19] ), 
            .\p[20] (\p[20] ), .\p[21] (\p[21] ), .\p[22] (\p[22] ), .\p[23] (\p[23] ), 
            .\p[24] (\p[24] ), .\p[25] (\p[25] ), .\p[26] (\p[26] ), .\p[27] (\p[27] ), 
            .\p[28] (\p[28] ), .\p[29] (\p[29] ), .\p[30] (\p[30] ), .\a[31] (\a[31] ), 
            .t({t}), .LM32D_DAT_O({LM32D_DAT_O}), .REF_CLK_c_enable_1221(REF_CLK_c_enable_1221), 
            .SHAREDBUS_DAT_O({SHAREDBUS_DAT_O}), .LM32D_SEL_O({LM32D_SEL_O}), 
            .\LM32D_ADR_O[0] (\LM32D_ADR_O[0] ), .\LM32D_CTI_O[0] (\LM32D_CTI_O[0] ), 
            .n38965(n38965), .LM32D_STB_O(LM32D_STB_O), .n21(n21), .\LM32D_ADR_O[1] (\LM32D_ADR_O[1] ), 
            .\LM32D_ADR_O[2] (\LM32D_ADR_O[2] ), .\next_cycle_type[2] (\next_cycle_type[2] ), 
            .\LM32D_ADR_O[4] (\LM32D_ADR_O[4] ), .\LM32D_ADR_O[5] (\LM32D_ADR_O[5] ), 
            .\d_adr_o_31__N_2278[5] (\d_adr_o_31__N_2278[5] ), .\LM32D_ADR_O[6] (\LM32D_ADR_O[6] ), 
            .\LM32D_ADR_O[7] (\LM32D_ADR_O[7] ), .\LM32D_ADR_O[8] (\LM32D_ADR_O[8] ), 
            .\LM32D_ADR_O[9] (\LM32D_ADR_O[9] ), .\d_adr_o_31__N_2278[9] (\d_adr_o_31__N_2278[9] ), 
            .\LM32D_ADR_O[10] (\LM32D_ADR_O[10] ), .\d_adr_o_31__N_2278[10] (\d_adr_o_31__N_2278[10] ), 
            .\LM32D_ADR_O[11] (\LM32D_ADR_O[11] ), .\LM32D_ADR_O[12] (\LM32D_ADR_O[12] ), 
            .\LM32D_ADR_O[13] (\LM32D_ADR_O[13] ), .\LM32D_ADR_O[14] (\LM32D_ADR_O[14] ), 
            .\LM32D_ADR_O[15] (\LM32D_ADR_O[15] ), .\LM32D_ADR_O[16] (\LM32D_ADR_O[16] ), 
            .\LM32D_ADR_O[17] (\LM32D_ADR_O[17] ), .\LM32D_ADR_O[18] (\LM32D_ADR_O[18] ), 
            .\LM32D_ADR_O[19] (\LM32D_ADR_O[19] ), .\LM32D_ADR_O[20] (\LM32D_ADR_O[20] ), 
            .\LM32D_ADR_O[21] (\LM32D_ADR_O[21] ), .\LM32D_ADR_O[22] (\LM32D_ADR_O[22] ), 
            .\LM32D_ADR_O[23] (\LM32D_ADR_O[23] ), .\LM32D_ADR_O[24] (\LM32D_ADR_O[24] ), 
            .\LM32D_ADR_O[25] (\LM32D_ADR_O[25] ), .\LM32D_ADR_O[26] (\LM32D_ADR_O[26] ), 
            .\LM32D_ADR_O[27] (\LM32D_ADR_O[27] ), .\LM32D_ADR_O[28] (\LM32D_ADR_O[28] ), 
            .\LM32D_ADR_O[29] (\LM32D_ADR_O[29] ), .\LM32D_ADR_O[30] (\LM32D_ADR_O[30] ), 
            .\LM32D_ADR_O[31] (\LM32D_ADR_O[31] ), .n41387(n41387), .n9(n9), 
            .\state[0] (\state[0] ), .\state[2] (\state[2] ), .flush_set({flush_set}), 
            .flush_set_8__N_2513({flush_set_8__N_2513}), .\dcache_refill_address[5] (\dcache_refill_address[5] ), 
            .\dcache_refill_address[9] (\dcache_refill_address[9] ), .\dcache_refill_address[10] (\dcache_refill_address[10] ), 
            .\tmem_write_address[1] (\tmem_write_address[1] ), .\tmem_write_address[5] (\tmem_write_address[5] ), 
            .\tmem_write_address[6] (\tmem_write_address[6] ), .\dmem_write_address[3] (\dmem_write_address[3] ), 
            .\dmem_write_address[7] (\dmem_write_address[7] ), .\dmem_write_address[8] (\dmem_write_address[8] ), 
            .jtag_reg_q({jtag_reg_q}), .jtag_reg_d({jtag_reg_d}), .REF_CLK_c_enable_1373(REF_CLK_c_enable_1373), 
            .n4626({n4626}), .rx_toggle_r_r(rx_toggle_r_r), .rx_toggle_r_r_r(rx_toggle_r_r_r), 
            .uart_tx_byte({uart_tx_byte}), .jrx_csr_read_data_8__N_3304(jrx_csr_read_data_8__N_3304), 
            .jtag_update_N_3371(jtag_update_N_3371), .\jtag_reg_addr_q[1] (jtag_reg_addr_q[1]), 
            .n30162(n30162), .n43(n43), .n29834(n29834), .n36337(n36337), 
            .SPI_INT_O_N_4422(SPI_INT_O_N_4422), .SPI_INT_O_N_4417(SPI_INT_O_N_4417), 
            .SPI_INT_O_N_4421(SPI_INT_O_N_4421), .\genblk1.wait_one_tick_done (\genblk1.wait_one_tick_done ), 
            .n6781(n6781), .n6764(n6764), .n6749(n6749), .n41410(n41410), 
            .n13990(n13990), .n32216(n32216), .\LM32I_CTI_O[0] (\LM32I_CTI_O[0] ), 
            .REF_CLK_c_enable_97(REF_CLK_c_enable_97), .n30900(n30900), 
            .pc_d({pc_d}), .REF_CLK_c_enable_1131(REF_CLK_c_enable_1131), 
            .n6760(n6760), .n45105(n45105), .n73(n73_adj_232), .n41461(n41461), 
            .\next_cycle_type[2]_adj_203 (\next_cycle_type[2]_adj_233 ), .n45080(n45080), 
            .n41390(n41390), .n5223(n5223), .n37955(n37955), .n37956(n37956), 
            .n37954(n37954), .n41345(n41345), .n41250(n41250), .n41251(n41251), 
            .n41279(n41279), .\LM32I_ADR_O[2] (\LM32I_ADR_O[2] ), .n45079(n45079), 
            .\reg_12[2] (\reg_12[2] ), .n2(n2), .\reg_12[12] (\reg_12[12] ), 
            .n40677(n40677), .\reg_12[29] (\reg_12[29] ), .n2_adj_204(n2_adj_234), 
            .\reg_12[3] (\reg_12[3] ), .n2_adj_205(n2_adj_235), .\reg_12[6] (\reg_12[6] ), 
            .n2_adj_206(n2_adj_236), .\reg_12[4] (\reg_12[4] ), .n2_adj_207(n2_adj_237), 
            .\reg_12[14] (\reg_12[14] ), .n2_adj_208(n2_adj_238), .n41429(n41429), 
            .\reg_12[22] (\reg_12[22] ), .n2_adj_209(n2_adj_239), .\reg_12[13] (\reg_12[13] ), 
            .n2_adj_210(n2_adj_240), .\reg_12[21] (\reg_12[21] ), .n2_adj_211(n2_adj_241), 
            .\reg_12[28] (\reg_12[28] ), .n2_adj_212(n2_adj_242), .\reg_12[11] (\reg_12[11] ), 
            .n2_adj_213(n2_adj_243), .\reg_12[18] (\reg_12[18] ), .n2_adj_214(n2_adj_244), 
            .\reg_12[25] (\reg_12[25] ), .n2_adj_215(n2_adj_245), .\reg_12[9] (\reg_12[9] ), 
            .n2_adj_216(n2_adj_246), .\reg_12[17] (\reg_12[17] ), .n2_adj_217(n2_adj_247), 
            .\reg_12[24] (\reg_12[24] ), .n2_adj_218(n2_adj_248), .\reg_12[7] (\reg_12[7] ), 
            .n2_adj_219(n2_adj_249), .\reg_12[15] (\reg_12[15] ), .n2_adj_220(n2_adj_250), 
            .n6589(n6589), .n6584(n6584), .n37179(n37179), .n6439(n6439), 
            .n6434(n6434), .n37177(n37177), .n6599(n6599), .n6594(n6594), 
            .n37180(n37180), .n6629(n6629), .n6624(n6624), .n37183(n37183), 
            .n6579(n6579), .n6574(n6574), .n37178(n37178), .n6429(n6429), 
            .n6424(n6424), .n37176(n37176), .n6609(n6609), .n6604(n6604), 
            .n37181(n37181), .n6619(n6619), .n6614(n6614), .n37182(n37182), 
            .n37185(n37185), .n37184(n37184), .n37188(n37188), .n37187(n37187), 
            .n37186(n37186), .n37189(n37189), .n7603(n7603), .n7571(n7571), 
            .n7607(n7607), .n7575(n7575), .n7606(n7606), .n7574(n7574), 
            .n7604(n7604), .n7572(n7572), .n7605(n7605), .n7573(n7573), 
            .n7608(n7608), .n7576(n7576), .n7602(n7602), .n7570(n7570), 
            .\selected_1__N_354[0] (\selected_1__N_354[0] ), .n7601(n7601), 
            .n7569(n7569), .n7600(n7600), .n7568(n7568), .n7599(n7599), 
            .n7567(n7567), .n7598(n7598), .n7566(n7566), .n7597(n7597), 
            .n7565(n7565), .n7596(n7596), .n7564(n7564), .n7595(n7595), 
            .n7563(n7563), .n7594(n7594), .n7562(n7562), .n7593(n7593), 
            .n7561(n7561), .n7592(n7592), .n7560(n7560), .n7584(n7584), 
            .n7552(n7552), .n7583(n7583), .n7551(n7551), .n7582(n7582), 
            .n7550(n7550), .n7581(n7581), .n7549(n7549), .n7580(n7580), 
            .n7548(n7548), .n7579(n7579), .n7547(n7547), .n7578(n7578), 
            .n7546(n7546), .n7577(n7577), .n7545(n7545), .n6750(n6750), 
            .n7591(n7591), .n7559(n7559), .n7590(n7590), .n7558(n7558), 
            .n7589(n7589), .n7557(n7557), .n7588(n7588), .n7556(n7556), 
            .n7587(n7587), .n7555(n7555), .n7586(n7586), .n7554(n7554), 
            .n7585(n7585), .n7553(n7553), .n37501(n37501), .n37500(n37500), 
            .n37502(n37502), .n37499(n37499), .n37498(n37498), .n37497(n37497), 
            .n37496(n37496), .n6751(n6751), .n6752(n6752), .n6753(n6753), 
            .n6754(n6754), .n6755(n6755), .n6756(n6756), .n6757(n6757), 
            .n6758(n6758), .n6759(n6759), .n6761(n6761), .n6762(n6762), 
            .n6763(n6763), .n37495(n37495), .n7672(n7672), .n7640(n7640), 
            .n7673(n7673), .n7641(n7641), .n34(n34), .n7674(n7674), 
            .n7642(n7642), .n7675(n7675), .n7643(n7643), .n7676(n7676), 
            .n7644(n7644), .n7671(n7671), .n7639(n7639), .n7670(n7670), 
            .n7638(n7638), .n7669(n7669), .n7637(n7637), .n7668(n7668), 
            .n7636(n7636), .n7667(n7667), .n7635(n7635), .n7666(n7666), 
            .n7634(n7634), .n7665(n7665), .n7633(n7633), .n7664(n7664), 
            .n7632(n7632), .n7663(n7663), .n7631(n7631), .n7662(n7662), 
            .n7630(n7630), .n7661(n7661), .n7629(n7629), .n7660(n7660), 
            .n7628(n7628), .n36(n36), .n7652(n7652), .n7620(n7620), 
            .n7651(n7651), .n7619(n7619), .n7650(n7650), .n7618(n7618), 
            .n7649(n7649), .n7617(n7617), .n37(n37), .n7648(n7648), 
            .n7616(n7616), .n7647(n7647), .n7615(n7615), .n7646(n7646), 
            .n7614(n7614), .n7645(n7645), .n7613(n7613), .n7659(n7659), 
            .n7627(n7627), .n7658(n7658), .n7626(n7626), .n7657(n7657), 
            .n7625(n7625), .n7656(n7656), .n7624(n7624), .n7655(n7655), 
            .n7623(n7623), .n7654(n7654), .n7622(n7622), .n7653(n7653), 
            .n7621(n7621), .n37504(n37504), .n37503(n37503), .n37507(n37507), 
            .n37506(n37506), .n37505(n37505), .n37508(n37508), .n45106(n45106), 
            .\LM32I_ADR_O[4] (\LM32I_ADR_O[4] ), .\LM32I_ADR_O[5] (\LM32I_ADR_O[5] ), 
            .\LM32I_ADR_O[6] (\LM32I_ADR_O[6] ), .\LM32I_ADR_O[7] (\LM32I_ADR_O[7] ), 
            .\LM32I_ADR_O[8] (\LM32I_ADR_O[8] ), .\LM32I_ADR_O[9] (\LM32I_ADR_O[9] ), 
            .\LM32I_ADR_O[10] (\LM32I_ADR_O[10] ), .\LM32I_ADR_O[11] (\LM32I_ADR_O[11] ), 
            .\LM32I_ADR_O[12] (\LM32I_ADR_O[12] ), .\LM32I_ADR_O[13] (\LM32I_ADR_O[13] ), 
            .\LM32I_ADR_O[14] (\LM32I_ADR_O[14] ), .\LM32I_ADR_O[15] (\LM32I_ADR_O[15] ), 
            .\LM32I_ADR_O[16] (\LM32I_ADR_O[16] ), .\LM32I_ADR_O[17] (\LM32I_ADR_O[17] ), 
            .\LM32I_ADR_O[18] (\LM32I_ADR_O[18] ), .\LM32I_ADR_O[19] (\LM32I_ADR_O[19] ), 
            .\LM32I_ADR_O[20] (\LM32I_ADR_O[20] ), .\LM32I_ADR_O[21] (\LM32I_ADR_O[21] ), 
            .\LM32I_ADR_O[22] (\LM32I_ADR_O[22] ), .\LM32I_ADR_O[23] (\LM32I_ADR_O[23] ), 
            .\LM32I_ADR_O[24] (\LM32I_ADR_O[24] ), .\LM32I_ADR_O[25] (\LM32I_ADR_O[25] ), 
            .\LM32I_ADR_O[26] (\LM32I_ADR_O[26] ), .\LM32I_ADR_O[27] (\LM32I_ADR_O[27] ), 
            .\LM32I_ADR_O[28] (\LM32I_ADR_O[28] ), .\LM32I_ADR_O[29] (\LM32I_ADR_O[29] ), 
            .\LM32I_ADR_O[30] (\LM32I_ADR_O[30] ), .\LM32I_ADR_O[31] (\LM32I_ADR_O[31] ), 
            .n949({n949}), .n32220(n32220), .selected({selected}), .flush_set_adj_231({flush_set_adj_272}), 
            .flush_set_8__N_1953({flush_set_8__N_1953}), .n157({n157}), 
            .n36336(n36336), .n10589(n10589), .n10585(n10585), .n10591(n10591), 
            .n10593(n10593), .n10587(n10587), .n10595(n10595), .n10452(n10452)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_top.v(283[10] 366[6])
    
endmodule
//
// Verilog Description of module jtag_cores
// module not written out since it is a black-box. 
//

//
// Verilog Description of module lm32_monitor
//

module lm32_monitor (REF_CLK_c, n69, ROM_ACK_O, REF_CLK_c_enable_1606, 
            state_1__N_3407, ROM_DAT_O, write_enable, n6362, n78, 
            n87, n96, \counter[2] , n41246, n19808, data, GND_net, 
            \SHAREDBUS_ADR_I[10] , n41310, n41301, \SHAREDBUS_ADR_I[7] , 
            n41346, \SHAREDBUS_ADR_I[5] , n41347, n41344, n41345, 
            VCC_net) /* synthesis syn_module_defined=1 */ ;
    input REF_CLK_c;
    input [7:0]n69;
    output ROM_ACK_O;
    input REF_CLK_c_enable_1606;
    output [1:0]state_1__N_3407;
    output [31:0]ROM_DAT_O;
    output write_enable;
    input n6362;
    input [7:0]n78;
    input [7:0]n87;
    input [7:0]n96;
    input \counter[2] ;
    input n41246;
    input n19808;
    output [31:0]data;
    input GND_net;
    input \SHAREDBUS_ADR_I[10] ;
    input n41310;
    input n41301;
    input \SHAREDBUS_ADR_I[7] ;
    input n41346;
    input \SHAREDBUS_ADR_I[5] ;
    input n41347;
    input n41344;
    input n41345;
    input VCC_net;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    wire [31:0]write_data;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(107[22:32])
    
    wire REF_CLK_c_enable_885;
    wire [1:0]state;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(104[11:16])
    wire [1:0]state_1__N_3407_c;
    
    wire REF_CLK_c_enable_1009, n6280;
    wire [31:0]n4034;
    
    wire REF_CLK_c_enable_917;
    
    FD1P3AX write_data_i0_i0 (.D(n69[0]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i0.GSR = "ENABLED";
    FD1S3DX MON_ACK_O_31 (.D(state_1__N_3407[1]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(ROM_ACK_O)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_ACK_O_31.GSR = "ENABLED";
    FD1S3DX state_i0 (.D(state_1__N_3407_c[0]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam state_i0.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i0 (.D(n4034[0]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i0.GSR = "ENABLED";
    FD1S3DX write_enable_30 (.D(n6362), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(write_enable)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_enable_30.GSR = "ENABLED";
    FD1P3AX write_data_i0_i1 (.D(n69[1]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i1.GSR = "ENABLED";
    FD1P3AX write_data_i0_i2 (.D(n69[2]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i2.GSR = "ENABLED";
    FD1P3AX write_data_i0_i3 (.D(n69[3]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i3.GSR = "ENABLED";
    FD1P3AX write_data_i0_i4 (.D(n69[4]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i4.GSR = "ENABLED";
    FD1P3AX write_data_i0_i5 (.D(n69[5]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i5.GSR = "ENABLED";
    FD1P3AX write_data_i0_i6 (.D(n69[6]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i6.GSR = "ENABLED";
    FD1P3AX write_data_i0_i7 (.D(n69[7]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i7.GSR = "ENABLED";
    FD1P3AX write_data_i0_i8 (.D(n78[0]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[8])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i8.GSR = "ENABLED";
    FD1P3AX write_data_i0_i9 (.D(n78[1]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[9])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i9.GSR = "ENABLED";
    FD1P3AX write_data_i0_i10 (.D(n78[2]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[10])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i10.GSR = "ENABLED";
    FD1P3AX write_data_i0_i11 (.D(n78[3]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[11])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i11.GSR = "ENABLED";
    FD1P3AX write_data_i0_i12 (.D(n78[4]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[12])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i12.GSR = "ENABLED";
    FD1P3AX write_data_i0_i13 (.D(n78[5]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[13])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i13.GSR = "ENABLED";
    FD1P3AX write_data_i0_i14 (.D(n78[6]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[14])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i14.GSR = "ENABLED";
    FD1P3AX write_data_i0_i15 (.D(n78[7]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[15])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i15.GSR = "ENABLED";
    FD1P3AX write_data_i0_i16 (.D(n87[0]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i16.GSR = "ENABLED";
    FD1P3AX write_data_i0_i17 (.D(n87[1]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i17.GSR = "ENABLED";
    FD1P3AX write_data_i0_i18 (.D(n87[2]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i18.GSR = "ENABLED";
    FD1P3AX write_data_i0_i19 (.D(n87[3]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i19.GSR = "ENABLED";
    FD1P3AX write_data_i0_i20 (.D(n87[4]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i20.GSR = "ENABLED";
    FD1P3AX write_data_i0_i21 (.D(n87[5]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i21.GSR = "ENABLED";
    FD1P3AX write_data_i0_i22 (.D(n87[6]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i22.GSR = "ENABLED";
    FD1P3AX write_data_i0_i23 (.D(n87[7]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i23.GSR = "ENABLED";
    FD1P3AX write_data_i0_i24 (.D(n96[0]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i24.GSR = "ENABLED";
    FD1P3AX write_data_i0_i25 (.D(n96[1]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i25.GSR = "ENABLED";
    FD1P3AX write_data_i0_i26 (.D(n96[2]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i26.GSR = "ENABLED";
    FD1P3AX write_data_i0_i27 (.D(n96[3]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i27.GSR = "ENABLED";
    FD1P3AX write_data_i0_i28 (.D(n96[4]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i28.GSR = "ENABLED";
    FD1P3AX write_data_i0_i29 (.D(n96[5]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i29.GSR = "ENABLED";
    FD1P3AX write_data_i0_i30 (.D(n96[6]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i30.GSR = "ENABLED";
    FD1P3AX write_data_i0_i31 (.D(n96[7]), .SP(REF_CLK_c_enable_885), .CK(REF_CLK_c), 
            .Q(write_data[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i31.GSR = "ENABLED";
    FD1P3DX state_i1 (.D(state_1__N_3407[1]), .SP(REF_CLK_c_enable_917), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam state_i1.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i1 (.D(n4034[1]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i1.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i2 (.D(n4034[2]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i2.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i3 (.D(n4034[3]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i3.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i4 (.D(n4034[4]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i4.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i5 (.D(n4034[5]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i5.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i6 (.D(n4034[6]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i6.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i7 (.D(n4034[7]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i7.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i8 (.D(n4034[8]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[8])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i8.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i9 (.D(n4034[9]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[9])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i9.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i10 (.D(n4034[10]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[10])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i10.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i11 (.D(n4034[11]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[11])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i11.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i12 (.D(n4034[12]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[12])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i12.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i13 (.D(n4034[13]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[13])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i13.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i14 (.D(n4034[14]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[14])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i14.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i15 (.D(n4034[15]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[15])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i15.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i16 (.D(n4034[16]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i16.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i17 (.D(n4034[17]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i17.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i18 (.D(n4034[18]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i18.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i19 (.D(n4034[19]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i19.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i20 (.D(n4034[20]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i20.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i21 (.D(n4034[21]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i21.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i22 (.D(n4034[22]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i22.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i23 (.D(n4034[23]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i23.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i24 (.D(n4034[24]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i24.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i25 (.D(n4034[25]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i25.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i26 (.D(n4034[26]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i26.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i27 (.D(n4034[27]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i27.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i28 (.D(n4034[28]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i28.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i29 (.D(n4034[29]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i29.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i30 (.D(n4034[30]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i30.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i31 (.D(n4034[31]), .SP(REF_CLK_c_enable_1009), .CD(n6280), 
            .CK(REF_CLK_c), .Q(ROM_DAT_O[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i31.GSR = "ENABLED";
    LUT4 i1_3_lut (.A(state[0]), .B(state[1]), .C(\counter[2] ), .Z(REF_CLK_c_enable_885)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut.init = 16'h2020;
    LUT4 i1_2_lut (.A(state[0]), .B(state[1]), .Z(state_1__N_3407[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam i1_2_lut.init = 16'h2222;
    LUT4 i12479_4_lut (.A(n41246), .B(state[1]), .C(state[0]), .D(n19808), 
         .Z(state_1__N_3407_c[0])) /* synthesis lut_function=(A (B (C)+!B !(C+(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(104[11:16])
    defparam i12479_4_lut.init = 16'hc0c2;
    LUT4 i14725_2_lut (.A(data[0]), .B(state[0]), .Z(n4034[0])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14725_2_lut.init = 16'h8888;
    LUT4 i33063_2_lut_rep_1004 (.A(state[0]), .B(state[1]), .Z(REF_CLK_c_enable_1009)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam i33063_2_lut_rep_1004.init = 16'h6666;
    LUT4 i1_3_lut_2_lut (.A(state[0]), .B(state[1]), .Z(n6280)) /* synthesis lut_function=(!(A+!(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam i1_3_lut_2_lut.init = 16'h4444;
    LUT4 i1_4_lut (.A(n41246), .B(state[1]), .C(n19808), .D(state[0]), 
         .Z(REF_CLK_c_enable_917)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B (D)+!B !(D)))) */ ;
    defparam i1_4_lut.init = 16'h3bce;
    LUT4 i14810_2_lut (.A(data[1]), .B(state[0]), .Z(n4034[1])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14810_2_lut.init = 16'h8888;
    LUT4 i14811_2_lut (.A(data[2]), .B(state[0]), .Z(n4034[2])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14811_2_lut.init = 16'h8888;
    LUT4 i14812_2_lut (.A(data[3]), .B(state[0]), .Z(n4034[3])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14812_2_lut.init = 16'h8888;
    LUT4 i14813_2_lut (.A(data[4]), .B(state[0]), .Z(n4034[4])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14813_2_lut.init = 16'h8888;
    LUT4 i14814_2_lut (.A(data[5]), .B(state[0]), .Z(n4034[5])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14814_2_lut.init = 16'h8888;
    LUT4 i14815_2_lut (.A(data[6]), .B(state[0]), .Z(n4034[6])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14815_2_lut.init = 16'h8888;
    LUT4 i14816_2_lut (.A(data[7]), .B(state[0]), .Z(n4034[7])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14816_2_lut.init = 16'h8888;
    LUT4 i14817_2_lut (.A(data[8]), .B(state[0]), .Z(n4034[8])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14817_2_lut.init = 16'h8888;
    LUT4 i14818_2_lut (.A(data[9]), .B(state[0]), .Z(n4034[9])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14818_2_lut.init = 16'h8888;
    LUT4 i14819_2_lut (.A(data[10]), .B(state[0]), .Z(n4034[10])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14819_2_lut.init = 16'h8888;
    LUT4 i14820_2_lut (.A(data[11]), .B(state[0]), .Z(n4034[11])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14820_2_lut.init = 16'h8888;
    LUT4 i14821_2_lut (.A(data[12]), .B(state[0]), .Z(n4034[12])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14821_2_lut.init = 16'h8888;
    LUT4 i14822_2_lut (.A(data[13]), .B(state[0]), .Z(n4034[13])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14822_2_lut.init = 16'h8888;
    LUT4 i14823_2_lut (.A(data[14]), .B(state[0]), .Z(n4034[14])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14823_2_lut.init = 16'h8888;
    LUT4 i14824_2_lut (.A(data[15]), .B(state[0]), .Z(n4034[15])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14824_2_lut.init = 16'h8888;
    LUT4 i14825_2_lut (.A(data[16]), .B(state[0]), .Z(n4034[16])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14825_2_lut.init = 16'h8888;
    LUT4 i14826_2_lut (.A(data[17]), .B(state[0]), .Z(n4034[17])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14826_2_lut.init = 16'h8888;
    LUT4 i14827_2_lut (.A(data[18]), .B(state[0]), .Z(n4034[18])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14827_2_lut.init = 16'h8888;
    LUT4 i14828_2_lut (.A(data[19]), .B(state[0]), .Z(n4034[19])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14828_2_lut.init = 16'h8888;
    LUT4 i14829_2_lut (.A(data[20]), .B(state[0]), .Z(n4034[20])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14829_2_lut.init = 16'h8888;
    LUT4 i14830_2_lut (.A(data[21]), .B(state[0]), .Z(n4034[21])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14830_2_lut.init = 16'h8888;
    LUT4 i14831_2_lut (.A(data[22]), .B(state[0]), .Z(n4034[22])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14831_2_lut.init = 16'h8888;
    LUT4 i14832_2_lut (.A(data[23]), .B(state[0]), .Z(n4034[23])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14832_2_lut.init = 16'h8888;
    LUT4 i14833_2_lut (.A(data[24]), .B(state[0]), .Z(n4034[24])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14833_2_lut.init = 16'h8888;
    LUT4 i14834_2_lut (.A(data[25]), .B(state[0]), .Z(n4034[25])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14834_2_lut.init = 16'h8888;
    LUT4 i14835_2_lut (.A(data[26]), .B(state[0]), .Z(n4034[26])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14835_2_lut.init = 16'h8888;
    LUT4 i14836_2_lut (.A(data[27]), .B(state[0]), .Z(n4034[27])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14836_2_lut.init = 16'h8888;
    LUT4 i14837_2_lut (.A(data[28]), .B(state[0]), .Z(n4034[28])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14837_2_lut.init = 16'h8888;
    LUT4 i14838_2_lut (.A(data[29]), .B(state[0]), .Z(n4034[29])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14838_2_lut.init = 16'h8888;
    LUT4 i14839_2_lut (.A(data[30]), .B(state[0]), .Z(n4034[30])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14839_2_lut.init = 16'h8888;
    LUT4 i14840_2_lut (.A(data[31]), .B(state[0]), .Z(n4034[31])) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i14840_2_lut.init = 16'h8888;
    lm32_monitor_ram ram (.write_data({write_data}), .GND_net(GND_net), 
            .\SHAREDBUS_ADR_I[10] (\SHAREDBUS_ADR_I[10] ), .n41310(n41310), 
            .n41301(n41301), .\SHAREDBUS_ADR_I[7] (\SHAREDBUS_ADR_I[7] ), 
            .n41346(n41346), .\SHAREDBUS_ADR_I[5] (\SHAREDBUS_ADR_I[5] ), 
            .n41347(n41347), .n41344(n41344), .n41345(n41345), .REF_CLK_c(REF_CLK_c), 
            .VCC_net(VCC_net), .write_enable(write_enable), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .data({data})) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(113[18] 130[6])
    
endmodule
//
// Verilog Description of module lm32_monitor_ram
//

module lm32_monitor_ram (write_data, GND_net, \SHAREDBUS_ADR_I[10] , n41310, 
            n41301, \SHAREDBUS_ADR_I[7] , n41346, \SHAREDBUS_ADR_I[5] , 
            n41347, n41344, n41345, REF_CLK_c, VCC_net, write_enable, 
            REF_CLK_c_enable_1606, data) /* synthesis syn_module_defined=1 */ ;
    input [31:0]write_data;
    input GND_net;
    input \SHAREDBUS_ADR_I[10] ;
    input n41310;
    input n41301;
    input \SHAREDBUS_ADR_I[7] ;
    input n41346;
    input \SHAREDBUS_ADR_I[5] ;
    input n41347;
    input n41344;
    input n41345;
    input REF_CLK_c;
    input VCC_net;
    input write_enable;
    input REF_CLK_c_enable_1606;
    output [31:0]data;
    
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    
    DP16KD \genblk1.lm32_monitor_ram_0_1_0  (.DIA0(write_data[18]), .DIA1(write_data[19]), 
           .DIA2(write_data[20]), .DIA3(write_data[21]), .DIA4(write_data[22]), 
           .DIA5(write_data[23]), .DIA6(write_data[24]), .DIA7(write_data[25]), 
           .DIA8(write_data[26]), .DIA9(write_data[27]), .DIA10(write_data[28]), 
           .DIA11(write_data[29]), .DIA12(write_data[30]), .DIA13(write_data[31]), 
           .DIA14(GND_net), .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), 
           .ADA0(VCC_net), .ADA1(VCC_net), .ADA2(GND_net), .ADA3(GND_net), 
           .ADA4(n41345), .ADA5(n41344), .ADA6(n41347), .ADA7(\SHAREDBUS_ADR_I[5] ), 
           .ADA8(n41346), .ADA9(\SHAREDBUS_ADR_I[7] ), .ADA10(n41301), 
           .ADA11(n41310), .ADA12(\SHAREDBUS_ADR_I[10] ), .ADA13(GND_net), 
           .CEA(VCC_net), .OCEA(VCC_net), .CLKA(REF_CLK_c), .WEA(write_enable), 
           .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), .RSTA(REF_CLK_c_enable_1606), 
           .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
           .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
           .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), 
           .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), 
           .DIB16(GND_net), .DIB17(GND_net), .ADB0(VCC_net), .ADB1(VCC_net), 
           .ADB2(GND_net), .ADB3(GND_net), .ADB4(GND_net), .ADB5(GND_net), 
           .ADB6(GND_net), .ADB7(GND_net), .ADB8(GND_net), .ADB9(GND_net), 
           .ADB10(GND_net), .ADB11(GND_net), .ADB12(GND_net), .ADB13(GND_net), 
           .CEB(GND_net), .OCEB(GND_net), .CLKB(REF_CLK_c), .WEB(GND_net), 
           .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), .RSTB(REF_CLK_c_enable_1606), 
           .DOA0(data[18]), .DOA1(data[19]), .DOA2(data[20]), .DOA3(data[21]), 
           .DOA4(data[22]), .DOA5(data[23]), .DOA6(data[24]), .DOA7(data[25]), 
           .DOA8(data[26]), .DOA9(data[27]), .DOA10(data[28]), .DOA11(data[29]), 
           .DOA12(data[30]), .DOA13(data[31])) /* synthesis MEM_LPC_FILE="lm32_monitor_ram.lpc", MEM_INIT_FILE="lm32_monitor.mem", syn_instantiated=1, LSE_LINE_FILE_ID=31, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=113, LSE_RLINE=130 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(113[18] 130[6])
    defparam \genblk1.lm32_monitor_ram_0_1_0 .DATA_WIDTH_A = 18;
    defparam \genblk1.lm32_monitor_ram_0_1_0 .DATA_WIDTH_B = 18;
    defparam \genblk1.lm32_monitor_ram_0_1_0 .REGMODE_A = "NOREG";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .REGMODE_B = "NOREG";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .RESETMODE = "SYNC";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .ASYNC_RESET_RELEASE = "SYNC";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .WRITEMODE_A = "NORMAL";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .WRITEMODE_B = "NORMAL";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .CSDECODE_A = "0b000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .CSDECODE_B = "0b000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .GSR = "ENABLED";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_00 = "0x0380003E0000D0802EE0016E703E0002EE80260000D0000D0000D0000D0000D0003E000340802600";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_01 = "0x0380003E0000D0802EE0016E703E0002EE8026000380003E0000D0802EE0016E703E0002EE802600";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_02 = "0x0380003E0000D0802EE0016E703E0002EE8026000380003E0000D0802EE0016E703E0002EE802600";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_03 = "0x0380003E0000D0802EE0016E703E0002EE8026000380003E0000D0802EE0016E703E0002EE802600";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_04 = "0x016EA016EA016E9016E9016E9016E9016E8016E8016E802600016E800DEF038FF00D0700DE702EE8";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_05 = "0x016EE016EE016ED016ED016ED016ED016EC016EC016EC016EC016EB016EB016EB016EB016EA016EA";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_06 = "0x00DE8016E802400016E802448016E802438016E802410016E802408016EF016EF016EF016EE016EE";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_07 = "0x00AE000AE000AE0030E800DEF02EE8016E8016E800AE8016E8000080000800008000080000800808";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_08 = "0x00AE400AE400AE400AE400AE300AE300AE300AE300AE200AE200AE200AE200AE100AE100AE100AE1";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_09 = "0x0340700AE70344F00AE70343F00AE700AE700AE700AE600AE600AE600AE600AE500AE500AE500AE5";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_0A = "0x00AE200AE200AE200AE200AE100AE100AE100AE100AE000AE000AE0030F000AE700AE70340F00AE7";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_0B = "0x00AE600AE600AE600AE600AE500AE500AE500AE500AE400AE400AE400AE400AE300AE300AE300AE3";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_0C = "0x011080081002478030F800AE700AE70340F00AE70340700AE70344F00AE70343F00AE700AE700AE7";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_0D = "0x016E700DE7030E8034700171002470030E80110801F0803470017100247000808030E80081003478";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_0E = "0x010E0016E0016E700DE7030E800DE700AE700AE000CE003EFF00CE003EFF00CE003EFF00CE003EFF";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_0F = "0x016E3016E3016E3016E3016E200DE7030E800DE700AE703EFF010E003EFF010E003EFF010E003EFF";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_10 = "0x00E7B01E0401E030347000D0001708024700347000D00017080247002E08016E7016E4016E4016E4";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_11 = "0x00D000170801F100110801F100110801F100110801F100110801F100110801F0802E0803EFF00E84";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_12 = "0x00AE400AE400AE400AE300AE300AE300AE300AE200D0000D0000D000342000D0000D0000D0003418";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_13 = "0x024500110C0287302430038FF03EFF02E700110801F100110801F0802E0803EFF030E800DE700AE7";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_14 = "0x0110801F100110801F100110801F100110801F100110801F0802E0803EFF02E0803EFF038FF02E70";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_15 = "0x03EFF02E88038FF034DA0170801F100110801F100110801F100110801F100110801F100110801F10";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_16 = "0x02E0803EFF02E0803EFF038FF00D5A03EFF00D63010580136300D0302E0803EFF02E0803EFF038FF";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_17 = "0x038FF0344A038FF03442038FF0343A038FF02E7002430038FF00D6300D5A00C5803EFF0136300D03";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_18 = "0x034D2038FF034C2038FF0349A038FF03EFF00D00038FF034CA038FF03492038FF0348A038FF03482";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_19 = "0x000000000000000000000000000000000000000000000000000000000000000000000000000038FF";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_0 .INIT_DATA = "STATIC";
    DP16KD \genblk1.lm32_monitor_ram_0_0_1  (.DIA0(write_data[0]), .DIA1(write_data[1]), 
           .DIA2(write_data[2]), .DIA3(write_data[3]), .DIA4(write_data[4]), 
           .DIA5(write_data[5]), .DIA6(write_data[6]), .DIA7(write_data[7]), 
           .DIA8(write_data[8]), .DIA9(write_data[9]), .DIA10(write_data[10]), 
           .DIA11(write_data[11]), .DIA12(write_data[12]), .DIA13(write_data[13]), 
           .DIA14(write_data[14]), .DIA15(write_data[15]), .DIA16(write_data[16]), 
           .DIA17(write_data[17]), .ADA0(VCC_net), .ADA1(VCC_net), .ADA2(GND_net), 
           .ADA3(GND_net), .ADA4(n41345), .ADA5(n41344), .ADA6(n41347), 
           .ADA7(\SHAREDBUS_ADR_I[5] ), .ADA8(n41346), .ADA9(\SHAREDBUS_ADR_I[7] ), 
           .ADA10(n41301), .ADA11(n41310), .ADA12(\SHAREDBUS_ADR_I[10] ), 
           .ADA13(GND_net), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(REF_CLK_c), 
           .WEA(write_enable), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(REF_CLK_c_enable_1606), .DIB0(GND_net), .DIB1(GND_net), 
           .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
           .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), 
           .DIB10(GND_net), .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), 
           .DIB14(GND_net), .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), 
           .ADB0(VCC_net), .ADB1(VCC_net), .ADB2(GND_net), .ADB3(GND_net), 
           .ADB4(GND_net), .ADB5(GND_net), .ADB6(GND_net), .ADB7(GND_net), 
           .ADB8(GND_net), .ADB9(GND_net), .ADB10(GND_net), .ADB11(GND_net), 
           .ADB12(GND_net), .ADB13(GND_net), .CEB(GND_net), .OCEB(GND_net), 
           .CLKB(REF_CLK_c), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
           .CSB2(GND_net), .RSTB(REF_CLK_c_enable_1606), .DOA0(data[0]), 
           .DOA1(data[1]), .DOA2(data[2]), .DOA3(data[3]), .DOA4(data[4]), 
           .DOA5(data[5]), .DOA6(data[6]), .DOA7(data[7]), .DOA8(data[8]), 
           .DOA9(data[9]), .DOA10(data[10]), .DOA11(data[11]), .DOA12(data[12]), 
           .DOA13(data[13]), .DOA14(data[14]), .DOA15(data[15]), .DOA16(data[16]), 
           .DOA17(data[17])) /* synthesis MEM_LPC_FILE="lm32_monitor_ram.lpc", MEM_INIT_FILE="lm32_monitor.mem", syn_instantiated=1, LSE_LINE_FILE_ID=31, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=113, LSE_RLINE=130 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(113[18] 130[6])
    defparam \genblk1.lm32_monitor_ram_0_0_1 .DATA_WIDTH_A = 18;
    defparam \genblk1.lm32_monitor_ram_0_0_1 .DATA_WIDTH_B = 18;
    defparam \genblk1.lm32_monitor_ram_0_0_1 .REGMODE_A = "NOREG";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .REGMODE_B = "NOREG";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .RESETMODE = "SYNC";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .ASYNC_RESET_RELEASE = "SYNC";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .WRITEMODE_A = "NORMAL";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .WRITEMODE_B = "NORMAL";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .CSDECODE_A = "0b000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .CSDECODE_B = "0b000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .GSR = "ENABLED";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_00 = "0x00096000EC1000400800300840003A000000000000000000000000000000000000003E0000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_01 = "0x00086000DC1000400800300840002A000000000000066000E4100040080020084000320000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_02 = "0x0004E000CC1000400800200840001A000000000000056000D4100040080020084000220000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_03 = "0x0003E000BC1000400800200840000A000000000000046000C4100040080020084000120000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_04 = "0x1002800024300202001C1001800014300102000C100080000000000106603FFC530000007F40E000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_05 = "0x1006800064300602005C1005800054300502004C1004800044300402003C1003800034300302002C";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_06 = "0x1F9A0100940080010090008001008C008001009C008001009800800300802007C00074300702006C";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_07 = "0x300102000C10008000001F9A00E000000041007810000100881000110001100011000110001100FF";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_08 = "0x300502004C1004800044300402003C1003800034300302002C1002800024300202001C1001800014";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_09 = "0x20000200942000020090200002008C3008010078300702006C1006800064300602005C1005800054";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_0A = "0x300302002C1002800024300202001C1001800014300102000C100080000000074200842000020098";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_0B = "0x300702006C1006800064300602005C1005800054300502004C1004800044300402003C1003800034";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_0C = "0x0FFFE1010001000000000007430084200002009830000300943000030090300003008C2007C10078";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_0D = "0x100040FFF400000200000FFFF01000000000000210054100000FFFF01000100FF00000100FF00000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_0E = "0x1000B10008100040FFF8000000000C1000410008100083FFE7100093FFE91000A3FFEB1000B3FFED";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_0F = "0x30014200181001C00020300240FFDC0000000008100043FFDD100083FFDF100093FFE11000A3FFE3";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_10 = "0x30000044003FC0010000100540FFFF0080010000100540FFFF008000880010004200081000C00010";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_11 = "0x100010FFF310063000501004D000471006D00046100720002C100570001F10077010003FFBC00000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_12 = "0x200081000C0001030014200181001C00020300240000000000000001000000000000000000010000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_13 = "0x070000FFFB30800070003FFD63FFB200800000041000A0004110006010003FF9A000000002410004";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_14 = "0x00033100110003310010000331000900033100080003310007010003FF89058003FF9C3FFF900800";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_15 = "0x3FF8D008003FFB4300000FFB61001B000361001A0002F10019000381001800038100130003310012";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_16 = "0x068003FF70058003FF723FFFB300013FF6A00001100001FFAB00000068003FF7B058003FF7D3FFB1";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_17 = "0x3FF92300003FF94300003FF96300003FFC100800070003FFFB0000130001100003FF5B1001700000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_18 = "0x300003FF83300003FF85300003FF873FF4A1004F3FF8A300003FF8C300003FF8E300003FF9030000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_19 = "0x0000000000000000000000000000000000000000000000000000000000000000000000000003FF81";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_1 .INIT_DATA = "STATIC";
    
endmodule
//
// Verilog Description of module lm32_cpu
//

module lm32_cpu (write_idx_w, n41352, n41351, w_result, n41350, REF_CLK_c, 
            REF_CLK_c_enable_1606, dcache_refill_request, \operand_1_x[1] , 
            dc_re, n41430, \counter[2] , n41432, REF_CLK_c_enable_176, 
            GND_net, n7611, n41405, REF_CLK_c_enable_164, n41380, 
            LM32D_CYC_O, locked_N_493, n41356, n41355, n41353, n41358, 
            n41359, \operand_m[10] , \operand_m[9] , \operand_m[5] , 
            LM32D_WE_O, dcache_select_x, n31750, n31955, n30241, n953, 
            n41326, n41354, bie, n31279, \adder_result_x[16] , \adder_result_x[17] , 
            \adder_result_x[18] , \adder_result_x[19] , \adder_result_x[20] , 
            \adder_result_x[21] , \adder_result_x[22] , \adder_result_x[23] , 
            \adder_result_x[24] , \adder_result_x[25] , \adder_result_x[26] , 
            \adder_result_x[27] , \adder_result_x[28] , \adder_result_x[29] , 
            \adder_result_x[30] , \adder_result_x[31] , n6518, n6648, 
            bus_error_f_N_1884, branch_target_d, direction_m, n45103, 
            n45099, n41394, n41401, bie_N_3274, pc_f, VCC_net, n41325, 
            n17816, n41379, \shifter_result_m[21] , \jtag_reg_addr_d[0] , 
            \jtag_reg_addr_d[1] , n41357, \left_shift_result[21] , \left_shift_result[10] , 
            b, \p[0] , \p[1] , \p[2] , \p[3] , \p[4] , \p[5] , 
            \p[6] , \p[7] , \p[8] , \p[9] , \p[10] , \p[11] , \p[12] , 
            \p[13] , \p[14] , \p[15] , \p[16] , \p[17] , \p[18] , 
            \p[19] , \p[20] , \p[21] , \p[22] , \p[23] , \p[24] , 
            \p[25] , \p[26] , \p[27] , \p[28] , \p[29] , \p[30] , 
            \a[31] , t, LM32D_DAT_O, REF_CLK_c_enable_1221, SHAREDBUS_DAT_O, 
            LM32D_SEL_O, \LM32D_ADR_O[0] , \LM32D_CTI_O[0] , n38965, 
            LM32D_STB_O, n21, \LM32D_ADR_O[1] , \LM32D_ADR_O[2] , \next_cycle_type[2] , 
            \LM32D_ADR_O[4] , \LM32D_ADR_O[5] , \d_adr_o_31__N_2278[5] , 
            \LM32D_ADR_O[6] , \LM32D_ADR_O[7] , \LM32D_ADR_O[8] , \LM32D_ADR_O[9] , 
            \d_adr_o_31__N_2278[9] , \LM32D_ADR_O[10] , \d_adr_o_31__N_2278[10] , 
            \LM32D_ADR_O[11] , \LM32D_ADR_O[12] , \LM32D_ADR_O[13] , \LM32D_ADR_O[14] , 
            \LM32D_ADR_O[15] , \LM32D_ADR_O[16] , \LM32D_ADR_O[17] , \LM32D_ADR_O[18] , 
            \LM32D_ADR_O[19] , \LM32D_ADR_O[20] , \LM32D_ADR_O[21] , \LM32D_ADR_O[22] , 
            \LM32D_ADR_O[23] , \LM32D_ADR_O[24] , \LM32D_ADR_O[25] , \LM32D_ADR_O[26] , 
            \LM32D_ADR_O[27] , \LM32D_ADR_O[28] , \LM32D_ADR_O[29] , \LM32D_ADR_O[30] , 
            \LM32D_ADR_O[31] , n41387, n9, \state[0] , \state[2] , 
            flush_set, flush_set_8__N_2513, \dcache_refill_address[5] , 
            \dcache_refill_address[9] , \dcache_refill_address[10] , \tmem_write_address[1] , 
            \tmem_write_address[5] , \tmem_write_address[6] , \dmem_write_address[3] , 
            \dmem_write_address[7] , \dmem_write_address[8] , jtag_reg_q, 
            jtag_reg_d, REF_CLK_c_enable_1373, n4626, rx_toggle_r_r, 
            rx_toggle_r_r_r, uart_tx_byte, jrx_csr_read_data_8__N_3304, 
            jtag_update_N_3371, \jtag_reg_addr_q[1] , n30162, n43, n29834, 
            n36337, SPI_INT_O_N_4422, SPI_INT_O_N_4417, SPI_INT_O_N_4421, 
            \genblk1.wait_one_tick_done , n6781, n6764, n6749, n41410, 
            n13990, n32216, \LM32I_CTI_O[0] , REF_CLK_c_enable_97, n30900, 
            pc_d, REF_CLK_c_enable_1131, n6760, n45105, n73, n41461, 
            \next_cycle_type[2]_adj_203 , n45080, n41390, n5223, n37955, 
            n37956, n37954, n41345, n41250, n41251, n41279, \LM32I_ADR_O[2] , 
            n45079, \reg_12[2] , n2, \reg_12[12] , n40677, \reg_12[29] , 
            n2_adj_204, \reg_12[3] , n2_adj_205, \reg_12[6] , n2_adj_206, 
            \reg_12[4] , n2_adj_207, \reg_12[14] , n2_adj_208, n41429, 
            \reg_12[22] , n2_adj_209, \reg_12[13] , n2_adj_210, \reg_12[21] , 
            n2_adj_211, \reg_12[28] , n2_adj_212, \reg_12[11] , n2_adj_213, 
            \reg_12[18] , n2_adj_214, \reg_12[25] , n2_adj_215, \reg_12[9] , 
            n2_adj_216, \reg_12[17] , n2_adj_217, \reg_12[24] , n2_adj_218, 
            \reg_12[7] , n2_adj_219, \reg_12[15] , n2_adj_220, n6589, 
            n6584, n37179, n6439, n6434, n37177, n6599, n6594, 
            n37180, n6629, n6624, n37183, n6579, n6574, n37178, 
            n6429, n6424, n37176, n6609, n6604, n37181, n6619, 
            n6614, n37182, n37185, n37184, n37188, n37187, n37186, 
            n37189, n7603, n7571, n7607, n7575, n7606, n7574, 
            n7604, n7572, n7605, n7573, n7608, n7576, n7602, n7570, 
            \selected_1__N_354[0] , n7601, n7569, n7600, n7568, n7599, 
            n7567, n7598, n7566, n7597, n7565, n7596, n7564, n7595, 
            n7563, n7594, n7562, n7593, n7561, n7592, n7560, n7584, 
            n7552, n7583, n7551, n7582, n7550, n7581, n7549, n7580, 
            n7548, n7579, n7547, n7578, n7546, n7577, n7545, n6750, 
            n7591, n7559, n7590, n7558, n7589, n7557, n7588, n7556, 
            n7587, n7555, n7586, n7554, n7585, n7553, n37501, 
            n37500, n37502, n37499, n37498, n37497, n37496, n6751, 
            n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, 
            n6761, n6762, n6763, n37495, n7672, n7640, n7673, 
            n7641, n34, n7674, n7642, n7675, n7643, n7676, n7644, 
            n7671, n7639, n7670, n7638, n7669, n7637, n7668, n7636, 
            n7667, n7635, n7666, n7634, n7665, n7633, n7664, n7632, 
            n7663, n7631, n7662, n7630, n7661, n7629, n7660, n7628, 
            n36, n7652, n7620, n7651, n7619, n7650, n7618, n7649, 
            n7617, n37, n7648, n7616, n7647, n7615, n7646, n7614, 
            n7645, n7613, n7659, n7627, n7658, n7626, n7657, n7625, 
            n7656, n7624, n7655, n7623, n7654, n7622, n7653, n7621, 
            n37504, n37503, n37507, n37506, n37505, n37508, n45106, 
            \LM32I_ADR_O[4] , \LM32I_ADR_O[5] , \LM32I_ADR_O[6] , \LM32I_ADR_O[7] , 
            \LM32I_ADR_O[8] , \LM32I_ADR_O[9] , \LM32I_ADR_O[10] , \LM32I_ADR_O[11] , 
            \LM32I_ADR_O[12] , \LM32I_ADR_O[13] , \LM32I_ADR_O[14] , \LM32I_ADR_O[15] , 
            \LM32I_ADR_O[16] , \LM32I_ADR_O[17] , \LM32I_ADR_O[18] , \LM32I_ADR_O[19] , 
            \LM32I_ADR_O[20] , \LM32I_ADR_O[21] , \LM32I_ADR_O[22] , \LM32I_ADR_O[23] , 
            \LM32I_ADR_O[24] , \LM32I_ADR_O[25] , \LM32I_ADR_O[26] , \LM32I_ADR_O[27] , 
            \LM32I_ADR_O[28] , \LM32I_ADR_O[29] , \LM32I_ADR_O[30] , \LM32I_ADR_O[31] , 
            n949, n32220, selected, flush_set_adj_231, flush_set_8__N_1953, 
            n157, n36336, n10589, n10585, n10591, n10593, n10587, 
            n10595, n10452) /* synthesis syn_module_defined=1 */ ;
    output [4:0]write_idx_w;
    output n41352;
    output n41351;
    output [31:0]w_result;
    output n41350;
    input REF_CLK_c;
    input REF_CLK_c_enable_1606;
    output dcache_refill_request;
    output \operand_1_x[1] ;
    output dc_re;
    output n41430;
    input \counter[2] ;
    input n41432;
    output REF_CLK_c_enable_176;
    input GND_net;
    output n7611;
    input n41405;
    output REF_CLK_c_enable_164;
    input n41380;
    output LM32D_CYC_O;
    output locked_N_493;
    output n41356;
    output n41355;
    output n41353;
    output n41358;
    output n41359;
    output \operand_m[10] ;
    output \operand_m[9] ;
    output \operand_m[5] ;
    output LM32D_WE_O;
    input dcache_select_x;
    input n31750;
    input n31955;
    input n30241;
    input [0:0]n953;
    input n41326;
    output n41354;
    output bie;
    output n31279;
    output \adder_result_x[16] ;
    output \adder_result_x[17] ;
    output \adder_result_x[18] ;
    output \adder_result_x[19] ;
    output \adder_result_x[20] ;
    output \adder_result_x[21] ;
    output \adder_result_x[22] ;
    output \adder_result_x[23] ;
    output \adder_result_x[24] ;
    output \adder_result_x[25] ;
    output \adder_result_x[26] ;
    output \adder_result_x[27] ;
    output \adder_result_x[28] ;
    output \adder_result_x[29] ;
    output \adder_result_x[30] ;
    output \adder_result_x[31] ;
    input n6518;
    input n6648;
    output bus_error_f_N_1884;
    input [31:2]branch_target_d;
    output direction_m;
    output n45103;
    output n45099;
    output n41394;
    output n41401;
    output bie_N_3274;
    output [31:2]pc_f;
    input VCC_net;
    output n41325;
    input n17816;
    output n41379;
    input \shifter_result_m[21] ;
    output \jtag_reg_addr_d[0] ;
    output \jtag_reg_addr_d[1] ;
    output n41357;
    output \left_shift_result[21] ;
    output \left_shift_result[10] ;
    output [31:0]b;
    output \p[0] ;
    output \p[1] ;
    output \p[2] ;
    output \p[3] ;
    output \p[4] ;
    output \p[5] ;
    output \p[6] ;
    output \p[7] ;
    output \p[8] ;
    output \p[9] ;
    output \p[10] ;
    output \p[11] ;
    output \p[12] ;
    output \p[13] ;
    output \p[14] ;
    output \p[15] ;
    output \p[16] ;
    output \p[17] ;
    output \p[18] ;
    output \p[19] ;
    output \p[20] ;
    output \p[21] ;
    output \p[22] ;
    output \p[23] ;
    output \p[24] ;
    output \p[25] ;
    output \p[26] ;
    output \p[27] ;
    output \p[28] ;
    output \p[29] ;
    output \p[30] ;
    output \a[31] ;
    input [32:0]t;
    output [31:0]LM32D_DAT_O;
    input REF_CLK_c_enable_1221;
    input [31:0]SHAREDBUS_DAT_O;
    output [3:0]LM32D_SEL_O;
    output \LM32D_ADR_O[0] ;
    output \LM32D_CTI_O[0] ;
    input n38965;
    output LM32D_STB_O;
    output n21;
    output \LM32D_ADR_O[1] ;
    output \LM32D_ADR_O[2] ;
    output \next_cycle_type[2] ;
    output \LM32D_ADR_O[4] ;
    output \LM32D_ADR_O[5] ;
    input \d_adr_o_31__N_2278[5] ;
    output \LM32D_ADR_O[6] ;
    output \LM32D_ADR_O[7] ;
    output \LM32D_ADR_O[8] ;
    output \LM32D_ADR_O[9] ;
    input \d_adr_o_31__N_2278[9] ;
    output \LM32D_ADR_O[10] ;
    input \d_adr_o_31__N_2278[10] ;
    output \LM32D_ADR_O[11] ;
    output \LM32D_ADR_O[12] ;
    output \LM32D_ADR_O[13] ;
    output \LM32D_ADR_O[14] ;
    output \LM32D_ADR_O[15] ;
    output \LM32D_ADR_O[16] ;
    output \LM32D_ADR_O[17] ;
    output \LM32D_ADR_O[18] ;
    output \LM32D_ADR_O[19] ;
    output \LM32D_ADR_O[20] ;
    output \LM32D_ADR_O[21] ;
    output \LM32D_ADR_O[22] ;
    output \LM32D_ADR_O[23] ;
    output \LM32D_ADR_O[24] ;
    output \LM32D_ADR_O[25] ;
    output \LM32D_ADR_O[26] ;
    output \LM32D_ADR_O[27] ;
    output \LM32D_ADR_O[28] ;
    output \LM32D_ADR_O[29] ;
    output \LM32D_ADR_O[30] ;
    output \LM32D_ADR_O[31] ;
    output n41387;
    input n9;
    output \state[0] ;
    output \state[2] ;
    output [8:0]flush_set;
    input [8:0]flush_set_8__N_2513;
    output \dcache_refill_address[5] ;
    output \dcache_refill_address[9] ;
    output \dcache_refill_address[10] ;
    input \tmem_write_address[1] ;
    input \tmem_write_address[5] ;
    input \tmem_write_address[6] ;
    input \dmem_write_address[3] ;
    input \dmem_write_address[7] ;
    input \dmem_write_address[8] ;
    input [7:0]jtag_reg_q;
    output [7:0]jtag_reg_d;
    input REF_CLK_c_enable_1373;
    input [7:0]n4626;
    output rx_toggle_r_r;
    output rx_toggle_r_r_r;
    output [7:0]uart_tx_byte;
    input jrx_csr_read_data_8__N_3304;
    input jtag_update_N_3371;
    input \jtag_reg_addr_q[1] ;
    input n30162;
    input n43;
    input n29834;
    input n36337;
    input SPI_INT_O_N_4422;
    input SPI_INT_O_N_4417;
    input SPI_INT_O_N_4421;
    output \genblk1.wait_one_tick_done ;
    output n6781;
    output n6764;
    output n6749;
    output n41410;
    input n13990;
    input n32216;
    output \LM32I_CTI_O[0] ;
    input REF_CLK_c_enable_97;
    input n30900;
    output [31:2]pc_d;
    input REF_CLK_c_enable_1131;
    output n6760;
    output n45105;
    input n73;
    output n41461;
    output \next_cycle_type[2]_adj_203 ;
    input n45080;
    input n41390;
    input n5223;
    output n37955;
    output n37956;
    output n37954;
    input n41345;
    output n41250;
    output n41251;
    output n41279;
    output \LM32I_ADR_O[2] ;
    input n45079;
    input \reg_12[2] ;
    output n2;
    input \reg_12[12] ;
    output n40677;
    input \reg_12[29] ;
    output n2_adj_204;
    input \reg_12[3] ;
    output n2_adj_205;
    input \reg_12[6] ;
    output n2_adj_206;
    input \reg_12[4] ;
    output n2_adj_207;
    input \reg_12[14] ;
    output n2_adj_208;
    input n41429;
    input \reg_12[22] ;
    output n2_adj_209;
    input \reg_12[13] ;
    output n2_adj_210;
    input \reg_12[21] ;
    output n2_adj_211;
    input \reg_12[28] ;
    output n2_adj_212;
    input \reg_12[11] ;
    output n2_adj_213;
    input \reg_12[18] ;
    output n2_adj_214;
    input \reg_12[25] ;
    output n2_adj_215;
    input \reg_12[9] ;
    output n2_adj_216;
    input \reg_12[17] ;
    output n2_adj_217;
    input \reg_12[24] ;
    output n2_adj_218;
    input \reg_12[7] ;
    output n2_adj_219;
    input \reg_12[15] ;
    output n2_adj_220;
    input n6589;
    input n6584;
    output n37179;
    input n6439;
    input n6434;
    output n37177;
    input n6599;
    input n6594;
    output n37180;
    input n6629;
    input n6624;
    output n37183;
    input n6579;
    input n6574;
    output n37178;
    input n6429;
    input n6424;
    output n37176;
    input n6609;
    input n6604;
    output n37181;
    input n6619;
    input n6614;
    output n37182;
    input n37185;
    input n37184;
    output n37188;
    input n37187;
    input n37186;
    output n37189;
    input n7603;
    input n7571;
    input n7607;
    input n7575;
    input n7606;
    input n7574;
    input n7604;
    input n7572;
    input n7605;
    input n7573;
    input n7608;
    input n7576;
    input n7602;
    input n7570;
    output \selected_1__N_354[0] ;
    input n7601;
    input n7569;
    input n7600;
    input n7568;
    input n7599;
    input n7567;
    input n7598;
    input n7566;
    input n7597;
    input n7565;
    input n7596;
    input n7564;
    input n7595;
    input n7563;
    input n7594;
    input n7562;
    input n7593;
    input n7561;
    input n7592;
    input n7560;
    input n7584;
    input n7552;
    input n7583;
    input n7551;
    input n7582;
    input n7550;
    input n7581;
    input n7549;
    input n7580;
    input n7548;
    input n7579;
    input n7547;
    input n7578;
    input n7546;
    input n7577;
    input n7545;
    output n6750;
    input n7591;
    input n7559;
    input n7590;
    input n7558;
    input n7589;
    input n7557;
    input n7588;
    input n7556;
    input n7587;
    input n7555;
    input n7586;
    input n7554;
    input n7585;
    input n7553;
    output n37501;
    output n37500;
    output n37502;
    output n37499;
    output n37498;
    output n37497;
    output n37496;
    output n6751;
    output n6752;
    output n6753;
    output n6754;
    output n6755;
    output n6756;
    output n6757;
    output n6758;
    output n6759;
    output n6761;
    output n6762;
    output n6763;
    output n37495;
    input n7672;
    input n7640;
    input n7673;
    input n7641;
    output n34;
    input n7674;
    input n7642;
    input n7675;
    input n7643;
    input n7676;
    input n7644;
    input n7671;
    input n7639;
    input n7670;
    input n7638;
    input n7669;
    input n7637;
    input n7668;
    input n7636;
    input n7667;
    input n7635;
    input n7666;
    input n7634;
    input n7665;
    input n7633;
    input n7664;
    input n7632;
    input n7663;
    input n7631;
    input n7662;
    input n7630;
    input n7661;
    input n7629;
    input n7660;
    input n7628;
    output n36;
    input n7652;
    input n7620;
    input n7651;
    input n7619;
    input n7650;
    input n7618;
    input n7649;
    input n7617;
    output n37;
    input n7648;
    input n7616;
    input n7647;
    input n7615;
    input n7646;
    input n7614;
    input n7645;
    input n7613;
    input n7659;
    input n7627;
    input n7658;
    input n7626;
    input n7657;
    input n7625;
    input n7656;
    input n7624;
    input n7655;
    input n7623;
    input n7654;
    input n7622;
    input n7653;
    input n7621;
    input n37504;
    input n37503;
    output n37507;
    input n37506;
    input n37505;
    output n37508;
    output n45106;
    output \LM32I_ADR_O[4] ;
    output \LM32I_ADR_O[5] ;
    output \LM32I_ADR_O[6] ;
    output \LM32I_ADR_O[7] ;
    output \LM32I_ADR_O[8] ;
    output \LM32I_ADR_O[9] ;
    output \LM32I_ADR_O[10] ;
    output \LM32I_ADR_O[11] ;
    output \LM32I_ADR_O[12] ;
    output \LM32I_ADR_O[13] ;
    output \LM32I_ADR_O[14] ;
    output \LM32I_ADR_O[15] ;
    output \LM32I_ADR_O[16] ;
    output \LM32I_ADR_O[17] ;
    output \LM32I_ADR_O[18] ;
    output \LM32I_ADR_O[19] ;
    output \LM32I_ADR_O[20] ;
    output \LM32I_ADR_O[21] ;
    output \LM32I_ADR_O[22] ;
    output \LM32I_ADR_O[23] ;
    output \LM32I_ADR_O[24] ;
    output \LM32I_ADR_O[25] ;
    output \LM32I_ADR_O[26] ;
    output \LM32I_ADR_O[27] ;
    output \LM32I_ADR_O[28] ;
    output \LM32I_ADR_O[29] ;
    output \LM32I_ADR_O[30] ;
    output \LM32I_ADR_O[31] ;
    input [0:0]n949;
    input n32220;
    input [1:0]selected;
    output [8:0]flush_set_adj_231;
    input [8:0]flush_set_8__N_1953;
    input [29:0]n157;
    input n36336;
    output n10589;
    output n10585;
    output n10591;
    output n10593;
    output n10587;
    output n10595;
    output n10452;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    wire jtag_update_N_3371 /* synthesis is_inv_clock=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(203[14:23])
    
    wire n35687;
    wire [31:0]w_result_31__N_690;
    wire [31:0]load_data_w;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(679[23:34])
    
    wire w_result_sel_load_w, raw_x_0, raw_m_0, n37947, n41232, n41233;
    wire [3:0]state;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(192[26:31])
    
    wire n32618;
    wire [31:0]operand_m;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(526[22:31])
    
    wire REF_CLK_c_enable_1235;
    wire [31:0]x_result;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(519[22:30])
    wire [4:0]write_idx_x;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(474[25:36])
    
    wire REF_CLK_c_enable_1624;
    wire [4:0]write_idx_d;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(473[26:37])
    wire [31:0]operand_0_x;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(523[22:33])
    
    wire REF_CLK_c_enable_4;
    wire [31:0]d_result_0;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(517[22:32])
    wire [31:8]deba;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(732[28:32])
    
    wire deba_31__N_1118;
    wire [31:0]operand_1_x;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(524[22:33])
    
    wire n37951, n37953, n37949, n41777;
    wire [31:0]adder_result_x;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(559[23:37])
    
    wire x_result_sel_add_x, n37950, n36552, n37952, n37948, data_bus_error_exception, 
        n6373, x_result_sel_csr_x, x_result_sel_sext_x, n37152, n37160, 
        x_result_sel_mc_arith_x, n36975, n36983, n36963, n36971, n36950, 
        n36958, n36937, n36945, n41400, valid_x, branch_flushX_m, 
        n20581, n36924, n36932, n36911, n36919, n36898, n36906, 
        cycles_5__N_2934, n31655, n36885, n36893, n36872, n36880, 
        n36859, n36867, n36846, n36854, n36833, n36841, REF_CLK_c_enable_61;
    wire [31:0]d_result_1;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(518[22:32])
    
    wire n36820, n36828, n36807, n36815, n36794, n36802, n36781, 
        n36789, w_result_sel_mul_x, w_result_sel_mul_d, n41775, n41773, 
        n41776, n36768, n36776, n36678, n36686, n36665, n36673, 
        valid_f, valid_f_N_1250, valid_a, w_result_sel_mul_m, n12394, 
        REF_CLK_c_enable_83, valid_x_N_1285, n36652, n36660;
    wire [1:0]size_x;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(392[22:28])
    
    wire n41366;
    wire [31:0]store_operand_x;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(525[22:37])
    wire [31:0]bypass_data_1;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(544[22:35])
    
    wire n36639, n36647;
    wire [31:2]branch_target_x;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(410[20:35])
    wire [29:0]branch_target_x_31__N_1120;
    wire [4:0]csr_x;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(478[22:27])
    wire [31:2]branch_target_m;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(411[20:35])
    wire [29:0]branch_target_m_31__N_1167;
    wire [31:8]eba;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(730[28:31])
    
    wire eba_31__N_1111;
    wire [31:0]operand_w;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(527[22:31])
    wire [31:0]operand_w_31__N_850;
    wire [4:0]write_idx_m;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(475[25:36])
    
    wire w_result_sel_load_m, w_result_sel_mul_w, write_enable_w, write_enable_m, 
        debug_exception_w, debug_exception_m, non_debug_exception_w, non_debug_exception_m, 
        n41203, interlock_N_1351, n30850, n12, n15;
    wire [31:2]memop_pc_w;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(514[20:30])
    
    wire memop_pc_w_31__N_1229;
    wire [31:2]pc_m;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(634[21:25])
    wire [4:0]write_idx_m_4__N_1162;
    
    wire valid_w, n30089, n32006, raw_x_1, load_d, n36627, n36635, 
        n36615, n36623, n31984, n31982, n36372, n36383, n32408, 
        n31831, n32404, n5915, n7;
    wire [31:0]n1261;
    
    wire n30245, n5, n31976, n41282, n22, REF_CLK_c_enable_712, 
        n36757, break_d, scall_d, n32142, eret_d, REF_CLK_c_enable_713, 
        n36746, csr_write_enable_x, n45068, n4, REF_CLK_c_enable_714, 
        w_result_sel_load_x, store_x, n36735, bret_d, bus_error_d, 
        n30070, REF_CLK_c_enable_715, n36724, n41499, n36713, REF_CLK_c_enable_460, 
        n36702, x_bypass_enable_x, x_bypass_enable_d, REF_CLK_c_enable_459, 
        n36691;
    wire [31:0]sext_result_x;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(572[23:36])
    wire [31:0]n5848;
    
    wire n27365, cmp_zero, dflush_m, n31501, n45171, REF_CLK_c_enable_1236, 
        valid_m, n30012, n3, n41575, n41572, n27364;
    wire [31:0]shifter_result_m;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(583[23:39])
    
    wire m_result_sel_shift_m, n41302, n27363, n35671, n32342, n2_c, 
        m_bypass_enable_x, m_bypass_enable_d, m_result_sel_shift_x;
    wire [31:0]n5814;
    wire [31:0]n5780;
    
    wire n40689, n40684;
    wire [2:0]condition_x;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(480[27:38])
    
    wire condition_met_x, n40686, n40685, n40687, n32262, n30479, 
        n4_adj_6193, n32258, n41731, n41727, n41732, reset_exception, 
        n12392, data_bus_error_exception_m, scall_x, n32260, branch_x, 
        branch_d, write_enable_x, write_enable_d, n35860, n2_adj_6194, 
        n32116, n35751, branch_taken_m_N_1388, exception_m, n30085, 
        branch_taken_m, adder_op_x, n41175, adder_op_x_n, adder_op_d_N_1366, 
        break_x, branch_predict_m, branch_predict_x, branch_predict_taken_m, 
        branch_predict_taken_x, load_m, store_m, write_enable_m_N_1339, 
        n41417, non_debug_exception_x, direction_x, n41365, store_d, 
        x_result_sel_csr_d, condition_met_m, n41184, branch_predict_taken_d, 
        m_result_sel_compare_x, m_result_sel_compare_d, eret_x, bret_x, 
        bus_error_x, eret_q_x, m_result_sel_shift_d, n41205, m_bypass_enable_m, 
        branch_m, m_result_sel_compare_m, REF_CLK_c_enable_430, REF_CLK_c_enable_431, 
        REF_CLK_c_enable_432, REF_CLK_c_enable_433, REF_CLK_c_enable_434, 
        REF_CLK_c_enable_435, REF_CLK_c_enable_436, REF_CLK_c_enable_437, 
        REF_CLK_c_enable_438, REF_CLK_c_enable_439, REF_CLK_c_enable_440, 
        REF_CLK_c_enable_441, REF_CLK_c_enable_442, REF_CLK_c_enable_443, 
        REF_CLK_c_enable_444, REF_CLK_c_enable_445, REF_CLK_c_enable_446, 
        REF_CLK_c_enable_447, REF_CLK_c_enable_448, REF_CLK_c_enable_449, 
        REF_CLK_c_enable_450, REF_CLK_c_enable_451, REF_CLK_c_enable_452, 
        REF_CLK_c_enable_453, REF_CLK_c_enable_454, REF_CLK_c_enable_388, 
        REF_CLK_c_enable_455, REF_CLK_c_enable_456, REF_CLK_c_enable_457, 
        REF_CLK_c_enable_458, n41295, n31334, REF_CLK_c_enable_1050, 
        n41231, n41197, REF_CLK_c_enable_1042, n30493, n7_adj_6195, 
        n41420, n12400, n11807, n35032, n35745, REF_CLK_c_enable_699, 
        REF_CLK_c_enable_700, REF_CLK_c_enable_701, REF_CLK_c_enable_702, 
        REF_CLK_c_enable_703, REF_CLK_c_enable_704, REF_CLK_c_enable_705, 
        REF_CLK_c_enable_706, REF_CLK_c_enable_707, REF_CLK_c_enable_708, 
        REF_CLK_c_enable_709, REF_CLK_c_enable_710, REF_CLK_c_enable_711, 
        REF_CLK_c_enable_716, REF_CLK_c_enable_717, REF_CLK_c_enable_718, 
        REF_CLK_c_enable_719, REF_CLK_c_enable_720, REF_CLK_c_enable_721, 
        REF_CLK_c_enable_722, REF_CLK_c_enable_723, REF_CLK_c_enable_724, 
        REF_CLK_c_enable_725, REF_CLK_c_enable_726, REF_CLK_c_enable_727, 
        REF_CLK_c_enable_728, REF_CLK_c_enable_729, n41367, data_bus_error_exception_N_1236, 
        n33176;
    wire [31:0]multiplier_result_w;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(597[23:42])
    
    wire n41391, n41240;
    wire [31:0]n4323;
    wire [31:0]ip;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(140[22:24])
    
    wire n41444;
    wire [31:0]x_result_31__N_1076;
    
    wire n36199;
    wire [31:0]x_result_31__N_626;
    
    wire n36268, n36247, n36196, n36223, n36283, n36244, n36184, 
        n36232, n36178, n36235, n36259, n36256, n36193, n36226, 
        n36187, n8, n36241, n36265, n36250, n36190, n36229, n36175, 
        n36238, n36262, n36253, REF_CLK_c_enable_823, REF_CLK_c_enable_1030, 
        n17970, n17971, n37174, n17972, n31825;
    wire [31:0]im;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(141[22:24])
    
    wire n41288, n31494, n12412, n12410, branch_flushX_m_N_1312, n31804, 
        n41450;
    wire [1:0]size_w;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(240[22:28])
    wire [31:0]data_w;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(248[22:28])
    
    wire n41164, n41160, n41156, n41152, n41148, n41144, n41140, 
        n41136, n41730, n41728, n41502, n41501, n41505, n41504, 
        n41508, n41507, n41511, n41510, n41168, n41514, n45175, 
        n35639, n41513, n41517, n41516;
    wire [2:0]state_adj_6256;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(186[26:31])
    
    wire n41520, n41519, n41523, n41522, n41526, n41525, n41529, 
        n41528, n41737, n41735, n41738, n41532, n41531, REF_CLK_c_enable_1299, 
        n41535, n41534, n41538, n41537, n41739, n41541, n41540, 
        n39321, n39320, n41741, n41544, stall_a, n41543, n41742;
    wire [10:0]\genblk1.ra ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(285[31:33])
    wire [10:0]n7388;
    
    wire n34890, n41547, n41546, n41743, n41550, n41549, n41553, 
        n41552, n7206;
    wire [10:0]n7190;
    
    wire n39330, n41556, n41555, n41744, n41745, n41559, n41558, 
        n7344;
    wire [10:0]n7322;
    
    wire n41562, n41561, n41565, n41564, n41746, n41568, n41567, 
        n39324, n39323, n41748, n7276;
    wire [10:0]n7256;
    wire [31:0]jrx_csr_read_data;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(686[23:40])
    
    wire n41571, n7274, n7272, n7270, n7220, n41308, n41570, n7356, 
        n41749, n7354, n7352, n41574, n41573, n41750, n7350, n41196, 
        n45181, n7348, REF_CLK_c_enable_1178, n7346, n7342, n45183, 
        n41138;
    wire [31:0]m_result;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(520[22:30])
    wire [31:0]bypass_data_0_31__N_882;
    
    wire n41283, n41217, REF_CLK_c_enable_1513;
    wire [31:0]n7609;
    
    wire raw_w_0;
    wire [31:0]bypass_data_0_31__N_1012;
    wire [31:0]bypass_data_1_31__N_914;
    wire [31:0]n7677;
    
    wire raw_w_1;
    wire [31:0]bypass_data_1_31__N_1044;
    
    wire n17969, n17974, n7338, stall_wb_load, n39333, n7340, n7336, 
        n7208, icache_refilling, dcache_refilling, n19852, n32128, 
        n32134, n32132, n33942, n33944, n33946, n7224, n41751, 
        n41752, n41142;
    wire [31:0]extended_immediate;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(324[23:41])
    
    wire n41179, n41375, n41291, n2_adj_6196, n41374, n2_adj_6197, 
        n41373, n2_adj_6198, n41372, n2_adj_6199, n41371, n2_adj_6200, 
        n41370, n2_adj_6201, n41361, n2_adj_6202, n41369, n2_adj_6203, 
        n41368, n2_adj_6204, n7222, n41348, n41198, n31335, n41377, 
        n2_adj_6205, n41376, n2_adj_6206, n7204, n7210, n7212, n7214, 
        n7216, n41388, n41389, n41215, REF_CLK_c_enable_1234;
    wire [31:0]bypass_data_0;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(543[22:35])
    
    wire n6026;
    wire [31:0]left_shift_result;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(93[22:39])
    
    wire n27362, n7218;
    wire [8:0]\genblk1.ra_adj_6257 ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(285[31:33])
    wire [8:0]n7502;
    
    wire n34898, n7290, n7288, n7286, n7284, n7282, n7280, n7278, 
        n32264, n41360, n9308, n41183, n41201, n32608, n19987, 
        n41146, valid_d, REF_CLK_c_enable_1622, n31132, n35022, n34986, 
        n35030, n41202;
    wire [31:0]dcache_refill_address;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(254[23:44])
    wire [31:0]d_adr_o_31__N_2278;
    
    wire n39310, n41150, n32630, n32636, n41216, n41435, n41154, 
        n41158, REF_CLK_c_enable_1425, n19, n41436, n17, n18, n41162, 
        n31549, n34880, REF_CLK_c_enable_1335, n41313, n34874, REF_CLK_c_enable_391, 
        n35412, n41753, n39327, n39326, n41755, ie, n9401, n41317, 
        jtag_reg_d_7__N_515, n41756, n41757, n41166, n41448, n41393, 
        n33932, n41758, n41759, n34936, n34942, n35767, n11934, 
        n27361, n41402, n27360, n27359, n41760, n39329, n41762, 
        n41763, n41764, n41208, n27358, n41765, n41766, n41413, 
        n34464, n41414, n41415, divide_by_zero_x;
    wire [2:0]eid_x_2__N_1009;
    
    wire n41772, jtag_break, n41767, n41774, n39332, REF_CLK_c_enable_1304;
    wire [31:0]logic_result_x;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(566[23:37])
    wire [2:0]eid_x_2__N_1108;
    
    wire n41416, n41498, n41284, adder_carry_n_x, n39318, n39317, 
        n41734, n41736;
    wire [31:0]operand_w_31__N_1197;
    
    wire n19316, n19330, n35587, n12404, n20639, REF_CLK_c_enable_949, 
        n41449, n41165, dcache_select_m, n30107, n41349, wb_select_m, 
        wb_load_complete, n41161, n19333, n19319, n41157, n41153, 
        n41729, n41149, n41145;
    wire [31:2]pc_x;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(633[21:25])
    wire [29:0]pc_a_31__N_1720;
    
    wire n41141, n31307, n37939, n31305, n31303, n2_adj_6216, n31301, 
        n2_adj_6217;
    wire [1:0]d_result_sel_1_d;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(413[33:49])
    
    wire n31299, n2_adj_6218, n31297, n2_adj_6219, n31324, n31312, 
        n31215, n37933, n31325, n31210, n31294, n31211, n37934, 
        n31308, n31209, n31318, n31207, n31314, n31214, n31296, 
        n31206, n37936, n31321, n37937, n31319, n31315, n31313, 
        n31311, n37938, n31295, n31306, n31317, n31320, n31309, 
        n31217, n31310, n31213, n31304, n31220, n37935, n31316, 
        n31212, n31302, n31216, n31322, n31221, n31300, n31219, 
        n31298, n31218, n31323, n31208, n41137, n37940, n37944, 
        n37946, n37942, n37943, n36614, n37945, n37941, n34556, 
        n2_adj_6220, n35591, raw_m_1, n35832, n33920, REF_CLK_c_enable_1366;
    wire [31:0]mc_result_x;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(616[23:34])
    
    wire q_d, n20863, n32652, n30879, icache_refill_request, dcache_restart_request, 
        icache_restart_request, n9304, n41187, n31996, way_match_0__N_2007, 
        n41178, n36389, n37914, n37915, n37919, n37917, n37916, 
        n37918, n41, restart_request_N_1998, n41172, n32278, n34542, 
        n6769, n45075, n41244, n41419, n41248, n30216, n6765, 
        n31717, n6771, n41228, n41437, n6778, n6780, n31542, n6768, 
        n32910, n6779, n10, n6777, n6775, n41382, n6770, n6766, 
        n6767, n6776, n40094, n41312, n41296, n41364, n41363, 
        n30820, n11834, n32356, n41281, n41441, n41229, n41227, 
        n41319, n41381, n41451, n41285, n30888, n41247;
    wire [31:0]instruction_d;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(654[30:43])
    
    wire n10475, n2_adj_6241, n2_adj_6242, n2_adj_6243, n2_adj_6244, 
        n6028, n40093, n10485, n31519, n30058, n41362, n41452, 
        n41241, n10_adj_6254, n41408;
    
    LUT4 i30528_4_lut (.A(write_idx_w[4]), .B(write_idx_w[2]), .C(n41352), 
         .D(n41351), .Z(n35687)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i30528_4_lut.init = 16'h7bde;
    PFUMX w_result_31__I_0_i4 (.BLUT(w_result_31__N_690[3]), .ALUT(load_data_w[3]), 
          .C0(w_result_sel_load_w), .Z(w_result[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i33184_rep_183_2_lut (.A(raw_x_0), .B(raw_m_0), .Z(n37947)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1516[10] 1521[36])
    defparam i33184_rep_183_2_lut.init = 16'heeee;
    LUT4 i1_3_lut_4_lut (.A(n41232), .B(n41233), .C(state[2]), .D(n41350), 
         .Z(n32618)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h2000;
    FD1P3DX operand_m_i0_i0 (.D(x_result[0]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i0.GSR = "ENABLED";
    FD1P3DX write_idx_x_i0_i0 (.D(write_idx_d[0]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(write_idx_x[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_x_i0_i0.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i0 (.D(d_result_0[0]), .SP(REF_CLK_c_enable_4), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i0.GSR = "ENABLED";
    FD1P3DX deba_i8_i8 (.D(operand_1_x[8]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[8])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i8.GSR = "ENABLED";
    LUT4 i33184_rep_187_2_lut (.A(raw_x_0), .B(raw_m_0), .Z(n37951)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1516[10] 1521[36])
    defparam i33184_rep_187_2_lut.init = 16'heeee;
    LUT4 i33184_rep_189_2_lut (.A(raw_x_0), .B(raw_m_0), .Z(n37953)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1516[10] 1521[36])
    defparam i33184_rep_189_2_lut.init = 16'heeee;
    LUT4 i33184_rep_185_2_lut (.A(raw_x_0), .B(raw_m_0), .Z(n37949)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1516[10] 1521[36])
    defparam i33184_rep_185_2_lut.init = 16'heeee;
    LUT4 n41777_bdd_3_lut (.A(n41777), .B(adder_result_x[14]), .C(x_result_sel_add_x), 
         .Z(x_result[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41777_bdd_3_lut.init = 16'hcaca;
    LUT4 i33184_rep_186_2_lut (.A(raw_x_0), .B(raw_m_0), .Z(n37950)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1516[10] 1521[36])
    defparam i33184_rep_186_2_lut.init = 16'heeee;
    LUT4 i33184_2_lut (.A(raw_x_0), .B(raw_m_0), .Z(n36552)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1516[10] 1521[36])
    defparam i33184_2_lut.init = 16'heeee;
    LUT4 i33184_rep_188_2_lut (.A(raw_x_0), .B(raw_m_0), .Z(n37952)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1516[10] 1521[36])
    defparam i33184_rep_188_2_lut.init = 16'heeee;
    LUT4 i33184_rep_184_2_lut (.A(raw_x_0), .B(raw_m_0), .Z(n37948)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1516[10] 1521[36])
    defparam i33184_rep_184_2_lut.init = 16'heeee;
    PFUMX w_result_31__I_0_i3 (.BLUT(w_result_31__N_690[2]), .ALUT(load_data_w[2]), 
          .C0(w_result_sel_load_w), .Z(w_result[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i2 (.BLUT(w_result_31__N_690[1]), .ALUT(load_data_w[1]), 
          .C0(w_result_sel_load_w), .Z(w_result[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1S3DX data_bus_error_seen_661 (.D(n6373), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(data_bus_error_exception)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2200[5] 2207[8])
    defparam data_bus_error_seen_661.GSR = "ENABLED";
    LUT4 i33284_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n37152), .Z(n37160)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(478[22:27])
    defparam i33284_4_lut.init = 16'hfffe;
    LUT4 i31980_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[3]), 
         .Z(n37152)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31980_2_lut.init = 16'h1111;
    LUT4 i33339_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36975), .Z(n36983)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33339_4_lut.init = 16'hfffe;
    LUT4 i31803_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[31]), 
         .Z(n36975)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31803_2_lut.init = 16'h1111;
    LUT4 i33341_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36963), .Z(n36971)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33341_4_lut.init = 16'hfffe;
    LUT4 i31791_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[30]), 
         .Z(n36963)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31791_2_lut.init = 16'h1111;
    LUT4 i33343_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36950), .Z(n36958)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33343_4_lut.init = 16'hfffe;
    LUT4 i31778_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[29]), 
         .Z(n36950)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31778_2_lut.init = 16'h1111;
    LUT4 i33345_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36937), .Z(n36945)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33345_4_lut.init = 16'hfffe;
    LUT4 i31765_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[28]), 
         .Z(n36937)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31765_2_lut.init = 16'h1111;
    LUT4 i1_2_lut_4_lut (.A(dcache_refill_request), .B(n41400), .C(valid_x), 
         .D(branch_flushX_m), .Z(n20581)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0040;
    LUT4 i33347_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36924), .Z(n36932)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33347_4_lut.init = 16'hfffe;
    LUT4 i31752_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[27]), 
         .Z(n36924)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31752_2_lut.init = 16'h1111;
    LUT4 i33349_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36911), .Z(n36919)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33349_4_lut.init = 16'hfffe;
    LUT4 i31739_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[26]), 
         .Z(n36911)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31739_2_lut.init = 16'h1111;
    LUT4 i33351_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36898), .Z(n36906)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33351_4_lut.init = 16'hfffe;
    LUT4 i31726_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[25]), 
         .Z(n36898)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31726_2_lut.init = 16'h1111;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(dcache_refill_request), .B(branch_flushX_m), 
         .C(valid_x), .D(cycles_5__N_2934), .Z(n31655)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'h1000;
    LUT4 i33353_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36885), .Z(n36893)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33353_4_lut.init = 16'hfffe;
    LUT4 i31713_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[24]), 
         .Z(n36885)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31713_2_lut.init = 16'h1111;
    LUT4 i33355_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36872), .Z(n36880)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33355_4_lut.init = 16'hfffe;
    LUT4 i31700_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[23]), 
         .Z(n36872)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31700_2_lut.init = 16'h1111;
    LUT4 i33357_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36859), .Z(n36867)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33357_4_lut.init = 16'hfffe;
    LUT4 i31687_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[22]), 
         .Z(n36859)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31687_2_lut.init = 16'h1111;
    LUT4 i33359_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36846), .Z(n36854)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33359_4_lut.init = 16'hfffe;
    LUT4 i31674_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[21]), 
         .Z(n36846)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31674_2_lut.init = 16'h1111;
    LUT4 i33361_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36833), .Z(n36841)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33361_4_lut.init = 16'hfffe;
    LUT4 i31661_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[20]), 
         .Z(n36833)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31661_2_lut.init = 16'h1111;
    FD1P3DX operand_1_x_i0_i0 (.D(d_result_1[0]), .SP(REF_CLK_c_enable_61), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i0.GSR = "ENABLED";
    LUT4 i33363_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36820), .Z(n36828)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33363_4_lut.init = 16'hfffe;
    LUT4 i31648_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[19]), 
         .Z(n36820)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31648_2_lut.init = 16'h1111;
    LUT4 i33365_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36807), .Z(n36815)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33365_4_lut.init = 16'hfffe;
    LUT4 i31635_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[18]), 
         .Z(n36807)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31635_2_lut.init = 16'h1111;
    LUT4 i33367_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36794), .Z(n36802)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33367_4_lut.init = 16'hfffe;
    LUT4 i31622_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[17]), 
         .Z(n36794)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31622_2_lut.init = 16'h1111;
    LUT4 i33369_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36781), .Z(n36789)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33369_4_lut.init = 16'hfffe;
    FD1P3DX w_result_sel_mul_x_679 (.D(w_result_sel_mul_d), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(w_result_sel_mul_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam w_result_sel_mul_x_679.GSR = "ENABLED";
    LUT4 i31609_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[16]), 
         .Z(n36781)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31609_2_lut.init = 16'h1111;
    LUT4 n41775_bdd_3_lut (.A(n41775), .B(n41773), .C(x_result_sel_sext_x), 
         .Z(n41776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41775_bdd_3_lut.init = 16'hcaca;
    LUT4 i33371_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36768), .Z(n36776)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33371_4_lut.init = 16'hfffe;
    LUT4 i31596_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[15]), 
         .Z(n36768)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31596_2_lut.init = 16'h1111;
    LUT4 i33088_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36678), .Z(n36686)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33088_4_lut.init = 16'hfffe;
    LUT4 i31506_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[7]), 
         .Z(n36678)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31506_2_lut.init = 16'h1111;
    LUT4 i33092_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36665), .Z(n36673)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33092_4_lut.init = 16'hfffe;
    LUT4 i31493_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[6]), 
         .Z(n36665)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31493_2_lut.init = 16'h1111;
    FD1P3DX valid_f_662 (.D(valid_a), .SP(valid_f_N_1250), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(valid_f)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2264[5] 2299[8])
    defparam valid_f_662.GSR = "ENABLED";
    FD1P3DX w_result_sel_mul_m_709 (.D(n12394), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(w_result_sel_mul_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam w_result_sel_mul_m_709.GSR = "ENABLED";
    FD1P3DX valid_x_664 (.D(valid_x_N_1285), .SP(REF_CLK_c_enable_83), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(valid_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2264[5] 2299[8])
    defparam valid_x_664.GSR = "ENABLED";
    LUT4 i33106_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36652), .Z(n36660)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33106_4_lut.init = 16'hfffe;
    LUT4 i31480_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[5]), 
         .Z(n36652)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31480_2_lut.init = 16'h1111;
    FD1P3DX size_x_i0_i0 (.D(n41366), .SP(REF_CLK_c_enable_1624), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(size_x[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam size_x_i0_i0.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i0 (.D(bypass_data_1[0]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i0.GSR = "ENABLED";
    LUT4 i33121_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36639), .Z(n36647)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33121_4_lut.init = 16'hfffe;
    FD1P3DX branch_target_x_i2_i2 (.D(branch_target_x_31__N_1120[0]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i2.GSR = "ENABLED";
    FD1P3DX csr_x_i0_i0 (.D(n41350), .SP(REF_CLK_c_enable_1624), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(csr_x[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam csr_x_i0_i0.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i2 (.D(branch_target_m_31__N_1167[0]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i2.GSR = "ENABLED";
    LUT4 i31467_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[4]), 
         .Z(n36639)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31467_2_lut.init = 16'h1111;
    FD1P3DX eba_i8_i8 (.D(operand_1_x[8]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[8])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i8.GSR = "ENABLED";
    FD1S3DX operand_w_i0 (.D(operand_w_31__N_850[0]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(operand_w[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i0.GSR = "ENABLED";
    FD1S3DX write_idx_w_i0 (.D(write_idx_m[0]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(write_idx_w[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_w_i0.GSR = "ENABLED";
    FD1S3DX w_result_sel_load_w_724 (.D(w_result_sel_load_m), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(w_result_sel_load_w)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam w_result_sel_load_w_724.GSR = "ENABLED";
    FD1S3DX w_result_sel_mul_w_725 (.D(w_result_sel_mul_m), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(w_result_sel_mul_w)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam w_result_sel_mul_w_725.GSR = "ENABLED";
    FD1S3DX write_enable_w_727 (.D(write_enable_m), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(write_enable_w)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_enable_w_727.GSR = "ENABLED";
    FD1S3DX debug_exception_w_728 (.D(debug_exception_m), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(debug_exception_w)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam debug_exception_w_728.GSR = "ENABLED";
    FD1S3DX non_debug_exception_w_729 (.D(non_debug_exception_m), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(non_debug_exception_w)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam non_debug_exception_w_729.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n41203), .B(interlock_N_1351), .C(n30850), .D(n12), 
         .Z(n15)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1873[20] 1904[21])
    defparam i1_4_lut.init = 16'h5554;
    FD1P3DX memop_pc_w_i2_i2 (.D(pc_m[2]), .SP(memop_pc_w_31__N_1229), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i2.GSR = "ENABLED";
    FD1P3DX write_idx_m_i0_i0 (.D(write_idx_m_4__N_1162[0]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(write_idx_m[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_m_i0_i0.GSR = "ENABLED";
    FD1S3DX valid_w_666 (.D(n30089), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(valid_w)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2264[5] 2299[8])
    defparam valid_w_666.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_584 (.A(n32006), .B(raw_x_1), .C(raw_x_0), .D(load_d), 
         .Z(interlock_N_1351)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1495[12] 1499[13])
    defparam i1_4_lut_adj_584.init = 16'ha0a8;
    LUT4 i33136_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36627), .Z(n36635)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33136_4_lut.init = 16'hfffe;
    LUT4 i31455_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[2]), 
         .Z(n36627)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31455_2_lut.init = 16'h1111;
    LUT4 i33149_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36615), .Z(n36623)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33149_4_lut.init = 16'hfffe;
    LUT4 i31443_2_lut (.A(x_result_sel_mc_arith_x), .B(\operand_1_x[1] ), 
         .Z(n36615)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31443_2_lut.init = 16'h1111;
    LUT4 i1_4_lut_adj_585 (.A(n31984), .B(n31982), .C(raw_m_0), .D(load_d), 
         .Z(n30850)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1501[16] 1503[17])
    defparam i1_4_lut_adj_585.init = 16'ha0a8;
    LUT4 i33236_4_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .D(n36372), .Z(n36383)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i33236_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_586 (.A(n32408), .B(n31831), .C(n32404), .D(branch_flushX_m), 
         .Z(n12)) /* synthesis lut_function=(A (B)+!A !(((D)+!C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1873[20] 1904[21])
    defparam i1_4_lut_adj_586.init = 16'h88c8;
    LUT4 i31200_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[0]), 
         .Z(n36372)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31200_2_lut.init = 16'h1111;
    LUT4 mux_75_i4_4_lut (.A(operand_0_x[3]), .B(n5915), .C(x_result_sel_csr_x), 
         .D(n7), .Z(n1261[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i4_4_lut.init = 16'hca0a;
    LUT4 i1_4_lut_adj_587 (.A(n30245), .B(n5), .C(n31976), .D(n41282), 
         .Z(n31982)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_587.init = 16'h0010;
    LUT4 i1_4_lut_adj_588 (.A(csr_x[4]), .B(n22), .C(csr_x[1]), .D(csr_x[2]), 
         .Z(n5915)) /* synthesis lut_function=(!(A+!(B (C (D))+!B (C+!(D))))) */ ;
    defparam i1_4_lut_adj_588.init = 16'h5011;
    LUT4 i27_3_lut (.A(csr_x[3]), .B(csr_x[1]), .C(csr_x[0]), .Z(n22)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_1115 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_712)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1115.init = 16'h0f0e;
    LUT4 i31585_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[14]), 
         .Z(n36757)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31585_2_lut.init = 16'h1111;
    LUT4 i1_4_lut_adj_589 (.A(break_d), .B(scall_d), .C(n32142), .D(eret_d), 
         .Z(n31831)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_589.init = 16'hfffe;
    LUT4 i1_2_lut_rep_1116 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_713)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1116.init = 16'h0f0e;
    LUT4 i31574_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[13]), 
         .Z(n36746)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31574_2_lut.init = 16'h1111;
    LUT4 i1_2_lut_3_lut (.A(csr_write_enable_x), .B(n45068), .C(csr_x[2]), 
         .Z(n4)) /* synthesis lut_function=(A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1983[31:78])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_1117 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_714)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1117.init = 16'h0f0e;
    LUT4 i1_4_lut_adj_590 (.A(dcache_refill_request), .B(w_result_sel_load_x), 
         .C(valid_x), .D(store_x), .Z(n32404)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;
    defparam i1_4_lut_adj_590.init = 16'h5040;
    LUT4 i31563_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[12]), 
         .Z(n36735)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31563_2_lut.init = 16'h1111;
    LUT4 i1_2_lut (.A(bret_d), .B(bus_error_d), .Z(n32142)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_591 (.A(dcache_refill_request), .B(branch_flushX_m), 
         .C(valid_x), .D(w_result_sel_load_x), .Z(n30070)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_591.init = 16'h1000;
    LUT4 i1_2_lut_rep_1118 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_715)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1118.init = 16'h0f0e;
    LUT4 i31552_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[11]), 
         .Z(n36724)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31552_2_lut.init = 16'h1111;
    LUT4 mux_508_i30_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[31]), .C(eba[31]), 
         .Z(n41499)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i30_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 i1_2_lut_rep_1119 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_4)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1119.init = 16'h0f0e;
    LUT4 i31541_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[10]), 
         .Z(n36713)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31541_2_lut.init = 16'h1111;
    LUT4 i1_2_lut_rep_1120 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_460)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1120.init = 16'h0f0e;
    LUT4 i31530_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[9]), 
         .Z(n36702)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31530_2_lut.init = 16'h1111;
    FD1P3DX x_bypass_enable_x_680 (.D(x_bypass_enable_d), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(x_bypass_enable_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam x_bypass_enable_x_680.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_1121 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_459)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1121.init = 16'h0f0e;
    LUT4 i31519_2_lut (.A(x_result_sel_mc_arith_x), .B(operand_1_x[8]), 
         .Z(n36691)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam i31519_2_lut.init = 16'h1111;
    LUT4 mux_75_i32_4_lut (.A(sext_result_x[31]), .B(n5848[31]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[31])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i32_4_lut.init = 16'hca0a;
    LUT4 mux_75_i31_4_lut (.A(sext_result_x[31]), .B(n5848[30]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[30])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i31_4_lut.init = 16'hca0a;
    LUT4 mux_75_i30_4_lut (.A(sext_result_x[31]), .B(n5848[29]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[29])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i30_4_lut.init = 16'hca0a;
    LUT4 mux_75_i29_4_lut (.A(sext_result_x[31]), .B(n5848[28]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[28])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i29_4_lut.init = 16'hca0a;
    LUT4 mux_75_i28_4_lut (.A(sext_result_x[31]), .B(n5848[27]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[27])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i28_4_lut.init = 16'hca0a;
    LUT4 mux_75_i27_4_lut (.A(sext_result_x[31]), .B(n5848[26]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[26])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i27_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_4_lut_adj_592 (.A(n41430), .B(dcache_refill_request), 
         .C(\counter[2] ), .D(n41432), .Z(REF_CLK_c_enable_176)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2700[10] 2703[12])
    defparam i1_2_lut_4_lut_adj_592.init = 16'h0020;
    LUT4 mux_75_i26_4_lut (.A(sext_result_x[31]), .B(n5848[25]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[25])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i26_4_lut.init = 16'hca0a;
    LUT4 mux_75_i25_4_lut (.A(sext_result_x[31]), .B(n5848[24]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[24])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i25_4_lut.init = 16'hca0a;
    LUT4 mux_75_i24_4_lut (.A(sext_result_x[31]), .B(n5848[23]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[23])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i24_4_lut.init = 16'hca0a;
    CCU2C operand_0_x_31__I_0_32 (.A0(\operand_1_x[1] ), .B0(operand_0_x[1]), 
          .C0(operand_1_x[0]), .D0(operand_0_x[0]), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n27365), .S1(cmp_zero));
    defparam operand_0_x_31__I_0_32.INIT0 = 16'h9009;
    defparam operand_0_x_31__I_0_32.INIT1 = 16'h0000;
    defparam operand_0_x_31__I_0_32.INJECT1_0 = "YES";
    defparam operand_0_x_31__I_0_32.INJECT1_1 = "NO";
    LUT4 mux_75_i23_4_lut (.A(sext_result_x[31]), .B(n5848[22]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[22])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i23_4_lut.init = 16'hca0a;
    FD1P3DX dflush_m_720 (.D(n31501), .SP(REF_CLK_c_enable_1235), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(dflush_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam dflush_m_720.GSR = "ENABLED";
    LUT4 i3148_2_lut_4_lut (.A(n41430), .B(dcache_refill_request), .C(\counter[2] ), 
         .D(write_idx_w[4]), .Z(n7611)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2700[10] 2703[12])
    defparam i3148_2_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_rep_840_4_lut (.A(n41430), .B(dcache_refill_request), 
         .C(\counter[2] ), .D(n41405), .Z(REF_CLK_c_enable_164)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2700[10] 2703[12])
    defparam i1_2_lut_rep_840_4_lut.init = 16'h0020;
    LUT4 i7032_2_lut_3_lut_4_lut (.A(n41380), .B(LM32D_CYC_O), .C(n45171), 
         .D(locked_N_493), .Z(REF_CLK_c_enable_1236)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2202[13:53])
    defparam i7032_2_lut_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i1_2_lut_adj_593 (.A(valid_m), .B(write_enable_m), .Z(n30012)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_593.init = 16'h8888;
    LUT4 mux_75_i22_4_lut (.A(sext_result_x[31]), .B(n5848[21]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[21])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i22_4_lut.init = 16'hca0a;
    LUT4 mux_75_i21_4_lut (.A(sext_result_x[31]), .B(n5848[20]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[20])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i21_4_lut.init = 16'hca0a;
    LUT4 i25228_4_lut (.A(write_idx_m[3]), .B(write_idx_m[0]), .C(n41356), 
         .D(n41355), .Z(n30245)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i25228_4_lut.init = 16'h7bde;
    LUT4 mux_75_i20_4_lut (.A(sext_result_x[31]), .B(n5848[19]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[19])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i20_4_lut.init = 16'hca0a;
    LUT4 mux_75_i19_4_lut (.A(sext_result_x[31]), .B(n5848[18]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[18])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i19_4_lut.init = 16'hca0a;
    LUT4 mux_75_i18_4_lut (.A(sext_result_x[31]), .B(n5848[17]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i18_4_lut.init = 16'hca0a;
    LUT4 mux_75_i17_4_lut (.A(sext_result_x[31]), .B(n5848[16]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[16])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i17_4_lut.init = 16'hca0a;
    LUT4 mux_75_i16_4_lut (.A(sext_result_x[31]), .B(n5848[15]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[15])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i16_4_lut.init = 16'hca0a;
    LUT4 mux_75_i8_4_lut (.A(operand_0_x[7]), .B(n5915), .C(x_result_sel_csr_x), 
         .D(n3), .Z(n1261[7])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i8_4_lut.init = 16'hca0a;
    LUT4 mux_75_i7_4_lut (.A(operand_0_x[6]), .B(n5848[6]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i7_4_lut.init = 16'hca0a;
    LUT4 mux_75_i6_4_lut (.A(operand_0_x[5]), .B(n41575), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[5])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i6_4_lut.init = 16'hca0a;
    LUT4 mux_75_i5_4_lut (.A(operand_0_x[4]), .B(n41572), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i5_4_lut.init = 16'hca0a;
    LUT4 mux_75_i3_4_lut (.A(operand_0_x[2]), .B(n5848[2]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i3_4_lut.init = 16'hca0a;
    LUT4 mux_75_i2_4_lut (.A(operand_0_x[1]), .B(n5848[1]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i2_4_lut.init = 16'hca0a;
    LUT4 mux_75_i1_4_lut (.A(operand_0_x[0]), .B(n5848[0]), .C(x_result_sel_csr_x), 
         .D(n5915), .Z(n1261[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i1_4_lut.init = 16'hca0a;
    CCU2C operand_0_x_31__I_0_31 (.A0(operand_1_x[5]), .B0(operand_0_x[5]), 
          .C0(operand_1_x[4]), .D0(operand_0_x[4]), .A1(operand_1_x[3]), 
          .B1(operand_0_x[3]), .C1(operand_1_x[2]), .D1(operand_0_x[2]), 
          .CIN(n27364), .COUT(n27365));
    defparam operand_0_x_31__I_0_31.INIT0 = 16'h9009;
    defparam operand_0_x_31__I_0_31.INIT1 = 16'h9009;
    defparam operand_0_x_31__I_0_31.INJECT1_0 = "YES";
    defparam operand_0_x_31__I_0_31.INJECT1_1 = "YES";
    LUT4 operand_m_31__I_0_744_i2_3_lut_rep_897 (.A(operand_m[1]), .B(shifter_result_m[1]), 
         .C(m_result_sel_shift_m), .Z(n41302)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1629[18] 1631[27])
    defparam operand_m_31__I_0_744_i2_3_lut_rep_897.init = 16'hcaca;
    CCU2C operand_0_x_31__I_0_29 (.A0(operand_1_x[9]), .B0(operand_0_x[9]), 
          .C0(operand_1_x[8]), .D0(operand_0_x[8]), .A1(operand_1_x[7]), 
          .B1(operand_0_x[7]), .C1(operand_1_x[6]), .D1(operand_0_x[6]), 
          .CIN(n27363), .COUT(n27364));
    defparam operand_0_x_31__I_0_29.INIT0 = 16'h9009;
    defparam operand_0_x_31__I_0_29.INIT1 = 16'h9009;
    defparam operand_0_x_31__I_0_29.INJECT1_0 = "YES";
    defparam operand_0_x_31__I_0_29.INJECT1_1 = "YES";
    LUT4 i1_4_lut_adj_594 (.A(n35671), .B(n32342), .C(write_idx_m[0]), 
         .D(n41350), .Z(raw_m_0)) /* synthesis lut_function=(!(A+!(B (C (D)+!C !(D))))) */ ;
    defparam i1_4_lut_adj_594.init = 16'h4004;
    LUT4 i30512_4_lut (.A(write_idx_m[4]), .B(write_idx_m[2]), .C(n41352), 
         .D(n41351), .Z(n35671)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i30512_4_lut.init = 16'h7bde;
    LUT4 i1_4_lut_adj_595 (.A(n2_c), .B(write_idx_m[3]), .C(n30012), .D(n41353), 
         .Z(n32342)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !((D)+!C)))) */ ;
    defparam i1_4_lut_adj_595.init = 16'h4010;
    FD1P3DX m_bypass_enable_x_681 (.D(m_bypass_enable_d), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(m_bypass_enable_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam m_bypass_enable_x_681.GSR = "ENABLED";
    FD1P3DX m_result_sel_shift_m_707 (.D(m_result_sel_shift_x), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(m_result_sel_shift_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam m_result_sel_shift_m_707.GSR = "ENABLED";
    PFUMX mux_2227_i1 (.BLUT(n5814[0]), .ALUT(n5780[0]), .C0(csr_x[2]), 
          .Z(n5848[0]));
    PFUMX i34158 (.BLUT(n40689), .ALUT(n40684), .C0(condition_x[2]), .Z(condition_met_x));
    PFUMX i34156 (.BLUT(n40686), .ALUT(n40685), .C0(cmp_zero), .Z(n40687));
    LUT4 i1_4_lut_adj_596 (.A(n32262), .B(n30479), .C(n4_adj_6193), .D(n32258), 
         .Z(raw_x_1)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_596.init = 16'h0010;
    LUT4 i1_4_lut_adj_597 (.A(write_idx_x[3]), .B(write_idx_x[1]), .C(n41356), 
         .D(n41358), .Z(n32258)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_597.init = 16'h7bde;
    PFUMX w_result_31__I_0_i1 (.BLUT(w_result_31__N_690[0]), .ALUT(load_data_w[0]), 
          .C0(w_result_sel_load_w), .Z(w_result[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX i34505 (.BLUT(n41731), .ALUT(n41727), .C0(x_result_sel_csr_x), 
          .Z(n41732));
    LUT4 i14612_3_lut (.A(data_bus_error_exception), .B(reset_exception), 
         .C(n45171), .Z(n12392)) /* synthesis lut_function=(!((B (C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i14612_3_lut.init = 16'h2a2a;
    FD1P3DX data_bus_error_exception_m_702 (.D(n12392), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(data_bus_error_exception_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam data_bus_error_exception_m_702.GSR = "ENABLED";
    FD1P3DX scall_x_698 (.D(scall_d), .SP(REF_CLK_c_enable_1624), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(scall_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam scall_x_698.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_598 (.A(write_idx_x[2]), .B(write_idx_x[0]), .C(n41359), 
         .D(n41355), .Z(n32260)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_598.init = 16'h7bde;
    FD1P3DX branch_x_693 (.D(branch_d), .SP(REF_CLK_c_enable_1624), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(branch_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_x_693.GSR = "ENABLED";
    FD1P3DX write_enable_x_682 (.D(write_enable_d), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(write_enable_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_enable_x_682.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_599 (.A(n35860), .B(n30479), .C(n2_adj_6194), .D(n32116), 
         .Z(raw_x_0)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_599.init = 16'h0100;
    LUT4 i30591_4_lut (.A(write_idx_x[4]), .B(write_idx_x[2]), .C(n41352), 
         .D(n41351), .Z(n35751)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i30591_4_lut.init = 16'h7bde;
    LUT4 i1_2_lut_adj_600 (.A(valid_x), .B(write_enable_x), .Z(n4_adj_6193)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_600.init = 16'h8888;
    LUT4 stall_m_N_1151_I_0_rep_104_4_lut (.A(n45171), .B(branch_taken_m_N_1388), 
         .C(exception_m), .D(n30085), .Z(branch_taken_m)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1655[30] 1668[31])
    defparam stall_m_N_1151_I_0_rep_104_4_lut.init = 16'ha8a0;
    FD1P3DX adder_op_x_689 (.D(n41175), .SP(REF_CLK_c_enable_1624), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(adder_op_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam adder_op_x_689.GSR = "ENABLED";
    FD1P3DX adder_op_x_n_690 (.D(adder_op_d_N_1366), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(adder_op_x_n)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam adder_op_x_n_690.GSR = "ENABLED";
    FD1P3DX break_x_697 (.D(break_d), .SP(REF_CLK_c_enable_1624), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(break_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam break_x_697.GSR = "ENABLED";
    FD1P3DX branch_predict_m_712 (.D(branch_predict_x), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_predict_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_predict_m_712.GSR = "ENABLED";
    FD1P3DX branch_predict_taken_m_713 (.D(branch_predict_taken_x), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_predict_taken_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_predict_taken_m_713.GSR = "ENABLED";
    FD1P3DX load_m_715 (.D(w_result_sel_load_x), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(load_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam load_m_715.GSR = "ENABLED";
    FD1P3DX store_m_716 (.D(store_x), .SP(REF_CLK_c_enable_1235), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(store_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_m_716.GSR = "ENABLED";
    FD1P3DX write_enable_m_717 (.D(write_enable_m_N_1339), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(write_enable_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_enable_m_717.GSR = "ENABLED";
    FD1P3DX debug_exception_m_721 (.D(n41417), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(debug_exception_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam debug_exception_m_721.GSR = "ENABLED";
    FD1P3DX non_debug_exception_m_722 (.D(non_debug_exception_x), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(non_debug_exception_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam non_debug_exception_m_722.GSR = "ENABLED";
    FD1P3DX direction_x_692 (.D(n41365), .SP(REF_CLK_c_enable_1624), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(direction_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam direction_x_692.GSR = "ENABLED";
    FD1P3DX store_x_686 (.D(store_d), .SP(REF_CLK_c_enable_1624), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(store_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_x_686.GSR = "ENABLED";
    FD1P3DX x_result_sel_csr_x_671 (.D(x_result_sel_csr_d), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(x_result_sel_csr_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam x_result_sel_csr_x_671.GSR = "ENABLED";
    FD1P3DX condition_met_m_719 (.D(condition_met_x), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(condition_met_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam condition_met_m_719.GSR = "ENABLED";
    FD1P3DX branch_predict_x_694 (.D(n41184), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_predict_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_predict_x_694.GSR = "ENABLED";
    FD1P3DX branch_predict_taken_x_695 (.D(branch_predict_taken_d), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_predict_taken_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_predict_taken_x_695.GSR = "ENABLED";
    FD1P3DX m_result_sel_compare_x_676 (.D(m_result_sel_compare_d), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(m_result_sel_compare_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam m_result_sel_compare_x_676.GSR = "ENABLED";
    FD1P3DX eret_x_699 (.D(eret_d), .SP(REF_CLK_c_enable_1624), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eret_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam eret_x_699.GSR = "ENABLED";
    FD1P3DX bret_x_700 (.D(bret_d), .SP(REF_CLK_c_enable_1624), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(bret_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam bret_x_700.GSR = "ENABLED";
    FD1P3DX bus_error_x_701 (.D(bus_error_d), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(bus_error_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam bus_error_x_701.GSR = "ENABLED";
    LUT4 eret_x_I_0_2_lut_4_lut (.A(dcache_refill_request), .B(branch_flushX_m), 
         .C(valid_x), .D(eret_x), .Z(eret_q_x)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam eret_x_I_0_2_lut_4_lut.init = 16'h1000;
    FD1P3DX m_result_sel_shift_x_677 (.D(m_result_sel_shift_d), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(m_result_sel_shift_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam m_result_sel_shift_x_677.GSR = "ENABLED";
    FD1P3DX csr_write_enable_x_703 (.D(n41205), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(csr_write_enable_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam csr_write_enable_x_703.GSR = "ENABLED";
    FD1P3DX m_bypass_enable_m_710 (.D(m_bypass_enable_x), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(m_bypass_enable_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam m_bypass_enable_m_710.GSR = "ENABLED";
    FD1P3DX branch_m_711 (.D(branch_x), .SP(REF_CLK_c_enable_1235), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(branch_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_m_711.GSR = "ENABLED";
    FD1P3DX m_result_sel_compare_m_706 (.D(m_result_sel_compare_x), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(m_result_sel_compare_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam m_result_sel_compare_m_706.GSR = "ENABLED";
    FD1P3DX w_result_sel_load_x_678 (.D(load_d), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(w_result_sel_load_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam w_result_sel_load_x_678.GSR = "ENABLED";
    FD1P3DX deba_i8_i31 (.D(operand_1_x[31]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i31.GSR = "ENABLED";
    FD1P3DX deba_i8_i30 (.D(operand_1_x[30]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i30.GSR = "ENABLED";
    FD1P3DX deba_i8_i29 (.D(operand_1_x[29]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i29.GSR = "ENABLED";
    FD1P3DX deba_i8_i28 (.D(operand_1_x[28]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i28.GSR = "ENABLED";
    FD1P3DX deba_i8_i27 (.D(operand_1_x[27]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i27.GSR = "ENABLED";
    FD1P3DX deba_i8_i26 (.D(operand_1_x[26]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i26.GSR = "ENABLED";
    FD1P3DX deba_i8_i25 (.D(operand_1_x[25]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i25.GSR = "ENABLED";
    FD1P3DX deba_i8_i24 (.D(operand_1_x[24]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i24.GSR = "ENABLED";
    FD1P3DX deba_i8_i23 (.D(operand_1_x[23]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i23.GSR = "ENABLED";
    FD1P3DX deba_i8_i22 (.D(operand_1_x[22]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i22.GSR = "ENABLED";
    FD1P3DX deba_i8_i21 (.D(operand_1_x[21]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i21.GSR = "ENABLED";
    FD1P3DX deba_i8_i20 (.D(operand_1_x[20]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i20.GSR = "ENABLED";
    FD1P3DX deba_i8_i19 (.D(operand_1_x[19]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i19.GSR = "ENABLED";
    FD1P3DX deba_i8_i18 (.D(operand_1_x[18]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i18.GSR = "ENABLED";
    FD1P3DX deba_i8_i17 (.D(operand_1_x[17]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i17.GSR = "ENABLED";
    FD1P3DX deba_i8_i16 (.D(operand_1_x[16]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i16.GSR = "ENABLED";
    FD1P3DX deba_i8_i15 (.D(operand_1_x[15]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[15])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i15.GSR = "ENABLED";
    FD1P3DX deba_i8_i14 (.D(operand_1_x[14]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[14])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i14.GSR = "ENABLED";
    FD1P3DX deba_i8_i13 (.D(operand_1_x[13]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[13])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i13.GSR = "ENABLED";
    FD1P3DX deba_i8_i12 (.D(operand_1_x[12]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[12])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i12.GSR = "ENABLED";
    FD1P3DX deba_i8_i11 (.D(operand_1_x[11]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[11])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i11.GSR = "ENABLED";
    FD1P3DX deba_i8_i10 (.D(operand_1_x[10]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[10])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i10.GSR = "ENABLED";
    FD1P3DX deba_i8_i9 (.D(operand_1_x[9]), .SP(deba_31__N_1118), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(deba[9])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i9.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i31 (.D(d_result_0[31]), .SP(REF_CLK_c_enable_430), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i31.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i30 (.D(d_result_0[30]), .SP(REF_CLK_c_enable_431), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i30.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i29 (.D(d_result_0[29]), .SP(REF_CLK_c_enable_432), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i29.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i28 (.D(d_result_0[28]), .SP(REF_CLK_c_enable_433), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i28.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i27 (.D(d_result_0[27]), .SP(REF_CLK_c_enable_434), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i27.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i26 (.D(d_result_0[26]), .SP(REF_CLK_c_enable_435), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i26.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i25 (.D(d_result_0[25]), .SP(REF_CLK_c_enable_436), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i25.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i24 (.D(d_result_0[24]), .SP(REF_CLK_c_enable_437), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i24.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i23 (.D(d_result_0[23]), .SP(REF_CLK_c_enable_438), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i23.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i22 (.D(d_result_0[22]), .SP(REF_CLK_c_enable_439), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i22.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i21 (.D(d_result_0[21]), .SP(REF_CLK_c_enable_440), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i21.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i20 (.D(d_result_0[20]), .SP(REF_CLK_c_enable_441), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i20.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i19 (.D(d_result_0[19]), .SP(REF_CLK_c_enable_442), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i19.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i18 (.D(d_result_0[18]), .SP(REF_CLK_c_enable_443), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i18.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i17 (.D(d_result_0[17]), .SP(REF_CLK_c_enable_444), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i17.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i16 (.D(d_result_0[16]), .SP(REF_CLK_c_enable_445), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i16.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i15 (.D(d_result_0[15]), .SP(REF_CLK_c_enable_446), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[15])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i15.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i14 (.D(d_result_0[14]), .SP(REF_CLK_c_enable_447), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[14])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i14.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i13 (.D(d_result_0[13]), .SP(REF_CLK_c_enable_448), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[13])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i13.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i12 (.D(d_result_0[12]), .SP(REF_CLK_c_enable_449), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[12])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i12.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i11 (.D(d_result_0[11]), .SP(REF_CLK_c_enable_450), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[11])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i11.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i10 (.D(d_result_0[10]), .SP(REF_CLK_c_enable_451), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[10])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i10.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i9 (.D(d_result_0[9]), .SP(REF_CLK_c_enable_452), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[9])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i9.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i8 (.D(d_result_0[8]), .SP(REF_CLK_c_enable_453), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[8])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i8.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i7 (.D(d_result_0[7]), .SP(REF_CLK_c_enable_454), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i7.GSR = "ENABLED";
    LUT4 csr_write_enable_x_I_0_2_lut_rep_802_4_lut (.A(dcache_refill_request), 
         .B(branch_flushX_m), .C(valid_x), .D(csr_write_enable_x), .Z(REF_CLK_c_enable_388)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam csr_write_enable_x_I_0_2_lut_rep_802_4_lut.init = 16'h1000;
    FD1P3DX operand_0_x_i0_i6 (.D(d_result_0[6]), .SP(REF_CLK_c_enable_455), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i6.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i5 (.D(d_result_0[5]), .SP(REF_CLK_c_enable_456), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i5.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i4 (.D(d_result_0[4]), .SP(REF_CLK_c_enable_457), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i4.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i3 (.D(d_result_0[3]), .SP(REF_CLK_c_enable_458), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i3.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i2 (.D(d_result_0[2]), .SP(REF_CLK_c_enable_459), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i2.GSR = "ENABLED";
    FD1P3DX operand_0_x_i0_i1 (.D(d_result_0[1]), .SP(REF_CLK_c_enable_460), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_0_x[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_0_x_i0_i1.GSR = "ENABLED";
    FD1P3DX write_idx_x_i0_i4 (.D(write_idx_d[4]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(write_idx_x[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_x_i0_i4.GSR = "ENABLED";
    FD1P3DX write_idx_x_i0_i3 (.D(write_idx_d[3]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(write_idx_x[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_x_i0_i3.GSR = "ENABLED";
    FD1P3DX write_idx_x_i0_i2 (.D(write_idx_d[2]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(write_idx_x[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_x_i0_i2.GSR = "ENABLED";
    FD1P3DX write_idx_x_i0_i1 (.D(write_idx_d[1]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(write_idx_x[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_x_i0_i1.GSR = "ENABLED";
    FD1P3DX condition_x_i0_i2 (.D(n41295), .SP(REF_CLK_c_enable_1624), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(condition_x[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam condition_x_i0_i2.GSR = "ENABLED";
    LUT4 i15529_rep_98_2_lut_4_lut (.A(dcache_refill_request), .B(branch_flushX_m), 
         .C(valid_x), .D(n41400), .Z(n31334)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i15529_rep_98_2_lut_4_lut.init = 16'h1000;
    FD1P3DX operand_m_i0_i31 (.D(x_result[31]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i31.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i30 (.D(x_result[30]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i30.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i29 (.D(x_result[29]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i29.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i28 (.D(x_result[28]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i28.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i27 (.D(x_result[27]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i27.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i26 (.D(x_result[26]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i26.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i25 (.D(x_result[25]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i25.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i24 (.D(x_result[24]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i24.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i23 (.D(x_result[23]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i23.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i22 (.D(x_result[22]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i22.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i21 (.D(x_result[21]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i21.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i20 (.D(x_result[20]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i20.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i19 (.D(x_result[19]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i19.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i18 (.D(x_result[18]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i18.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i17 (.D(x_result[17]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i17.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i16 (.D(x_result[16]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i16.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i15 (.D(x_result[15]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[15])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i15.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i14 (.D(x_result[14]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[14])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i14.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i13 (.D(x_result[13]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[13])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i13.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i12 (.D(x_result[12]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[12])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i12.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i11 (.D(x_result[11]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[11])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i11.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i10 (.D(x_result[10]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\operand_m[10] )) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i10.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i9 (.D(x_result[9]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\operand_m[9] )) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i9.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i8 (.D(x_result[8]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[8])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i8.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i7 (.D(x_result[7]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i7.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i6 (.D(x_result[6]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i6.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i5 (.D(x_result[5]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\operand_m[5] )) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i5.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i4 (.D(x_result[4]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i4.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i3 (.D(x_result[3]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i3.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i2 (.D(x_result[2]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i2.GSR = "ENABLED";
    FD1P3DX operand_m_i0_i1 (.D(x_result[1]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_m[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i1.GSR = "ENABLED";
    LUT4 branch_flushX_m_I_0_774_2_lut_rep_826 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .Z(n41231)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam branch_flushX_m_I_0_774_2_lut_rep_826.init = 16'heeee;
    LUT4 stall_m_I_0_745_2_lut_rep_792_3_lut_4_lut (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(n41197)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam stall_m_I_0_745_2_lut_rep_792_3_lut_4_lut.init = 16'hf0f1;
    LUT4 i1_2_lut_rep_785_3_lut_4_lut (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_1042)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_785_3_lut_4_lut.init = 16'h0f0e;
    LUT4 i14584_rep_827 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(cycles_5__N_2934), .Z(n41232)) /* synthesis lut_function=(A+(B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i14584_rep_827.init = 16'hfefe;
    LUT4 i33171_3_lut_4_lut_4_lut (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(cycles_5__N_2934), .D(n41233), .Z(REF_CLK_c_enable_83)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i33171_3_lut_4_lut_4_lut.init = 16'heefe;
    LUT4 i14685_2_lut_4_lut (.A(n30493), .B(n7_adj_6195), .C(n41420), 
         .D(LM32D_WE_O), .Z(n12400)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B (C+(D))))) */ ;
    defparam i14685_2_lut_4_lut.init = 16'h00ef;
    LUT4 i1_2_lut_rep_1122 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_458)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1122.init = 16'h0f0e;
    LUT4 i1_2_lut_4_lut_adj_601 (.A(n30493), .B(n7_adj_6195), .C(n41420), 
         .D(n11807), .Z(n35032)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_2_lut_4_lut_adj_601.init = 16'hffef;
    LUT4 i30585_2_lut_4_lut (.A(n30493), .B(n7_adj_6195), .C(n41420), 
         .D(dcache_select_x), .Z(n35745)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i30585_2_lut_4_lut.init = 16'hffef;
    FD1P3DX operand_1_x_i0_i1 (.D(d_result_1[1]), .SP(REF_CLK_c_enable_699), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\operand_1_x[1] )) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i1.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i2 (.D(d_result_1[2]), .SP(REF_CLK_c_enable_700), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i2.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i3 (.D(d_result_1[3]), .SP(REF_CLK_c_enable_701), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i3.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i4 (.D(d_result_1[4]), .SP(REF_CLK_c_enable_702), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i4.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i5 (.D(d_result_1[5]), .SP(REF_CLK_c_enable_703), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i5.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i6 (.D(d_result_1[6]), .SP(REF_CLK_c_enable_704), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i6.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i7 (.D(d_result_1[7]), .SP(REF_CLK_c_enable_705), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i7.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i8 (.D(d_result_1[8]), .SP(REF_CLK_c_enable_706), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[8])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i8.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i9 (.D(d_result_1[9]), .SP(REF_CLK_c_enable_707), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[9])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i9.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i10 (.D(d_result_1[10]), .SP(REF_CLK_c_enable_708), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[10])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i10.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i11 (.D(d_result_1[11]), .SP(REF_CLK_c_enable_709), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[11])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i11.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i12 (.D(d_result_1[12]), .SP(REF_CLK_c_enable_710), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[12])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i12.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i13 (.D(d_result_1[13]), .SP(REF_CLK_c_enable_711), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[13])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i13.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i14 (.D(d_result_1[14]), .SP(REF_CLK_c_enable_712), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[14])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i14.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i15 (.D(d_result_1[15]), .SP(REF_CLK_c_enable_713), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[15])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i15.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i16 (.D(d_result_1[16]), .SP(REF_CLK_c_enable_714), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i16.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i17 (.D(d_result_1[17]), .SP(REF_CLK_c_enable_715), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i17.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i18 (.D(d_result_1[18]), .SP(REF_CLK_c_enable_716), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i18.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i19 (.D(d_result_1[19]), .SP(REF_CLK_c_enable_717), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i19.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i20 (.D(d_result_1[20]), .SP(REF_CLK_c_enable_718), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i20.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i21 (.D(d_result_1[21]), .SP(REF_CLK_c_enable_719), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i21.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i22 (.D(d_result_1[22]), .SP(REF_CLK_c_enable_720), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i22.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i23 (.D(d_result_1[23]), .SP(REF_CLK_c_enable_721), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i23.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i24 (.D(d_result_1[24]), .SP(REF_CLK_c_enable_722), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i24.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i25 (.D(d_result_1[25]), .SP(REF_CLK_c_enable_723), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i25.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i26 (.D(d_result_1[26]), .SP(REF_CLK_c_enable_724), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i26.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i27 (.D(d_result_1[27]), .SP(REF_CLK_c_enable_725), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i27.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i28 (.D(d_result_1[28]), .SP(REF_CLK_c_enable_726), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i28.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i29 (.D(d_result_1[29]), .SP(REF_CLK_c_enable_727), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i29.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i30 (.D(d_result_1[30]), .SP(REF_CLK_c_enable_728), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i30.GSR = "ENABLED";
    FD1P3DX operand_1_x_i0_i31 (.D(d_result_1[31]), .SP(REF_CLK_c_enable_729), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(operand_1_x[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i31.GSR = "ENABLED";
    FD1P3DX size_x_i0_i1 (.D(n41367), .SP(REF_CLK_c_enable_1624), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(size_x[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam size_x_i0_i1.GSR = "ENABLED";
    LUT4 i14564_4_lut (.A(data_bus_error_exception), .B(data_bus_error_exception_N_1236), 
         .C(n33176), .D(n31750), .Z(n6373)) /* synthesis lut_function=(!(A (B)+!A (B+((D)+!C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2200[5] 2207[8])
    defparam i14564_4_lut.init = 16'h2232;
    LUT4 exception_m_I_0_800_2_lut (.A(exception_m), .B(dcache_refill_request), 
         .Z(data_bus_error_exception_N_1236)) /* synthesis lut_function=(!((B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2205[13:57])
    defparam exception_m_I_0_800_2_lut.init = 16'h2222;
    LUT4 i1_4_lut_adj_602 (.A(n31955), .B(n30241), .C(n953[0]), .D(n41326), 
         .Z(n33176)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2202[13:53])
    defparam i1_4_lut_adj_602.init = 16'h4000;
    LUT4 operand_w_31__I_0_i4_3_lut (.A(operand_w[3]), .B(multiplier_result_w[3]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_1123 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_457)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1123.init = 16'h0f0e;
    LUT4 i15314_4_lut_4_lut (.A(n41391), .B(n41240), .C(n4323[1]), .D(ip[1]), 
         .Z(n5814[1])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i15314_4_lut_4_lut.init = 16'h5140;
    LUT4 i32776_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[7]), 
         .D(n36199), .Z(x_result_31__N_626[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32776_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32808_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[30]), 
         .D(n36268), .Z(x_result_31__N_626[30])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32808_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32794_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[23]), 
         .D(n36247), .Z(x_result_31__N_626[23])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32794_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32774_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[6]), 
         .D(n36196), .Z(x_result_31__N_626[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32774_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32778_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[15]), 
         .D(n36223), .Z(x_result_31__N_626[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32778_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32810_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[31]), 
         .D(n36283), .Z(x_result_31__N_626[31])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32810_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32792_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[22]), 
         .D(n36244), .Z(x_result_31__N_626[22])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32792_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32768_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[2]), 
         .D(n36184), .Z(x_result_31__N_626[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32768_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32784_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[18]), 
         .D(n36232), .Z(x_result_31__N_626[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32784_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32766_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[1]), 
         .D(n36178), .Z(x_result_31__N_626[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32766_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32786_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[19]), 
         .D(n36235), .Z(x_result_31__N_626[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32786_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32802_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[27]), 
         .D(n36259), .Z(x_result_31__N_626[27])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32802_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32800_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[26]), 
         .D(n36256), .Z(x_result_31__N_626[26])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32800_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32772_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[5]), 
         .D(n36193), .Z(x_result_31__N_626[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32772_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32780_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[16]), 
         .D(n36226), .Z(x_result_31__N_626[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32780_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32812_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[3]), 
         .D(n36187), .Z(n8)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32812_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32790_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[21]), 
         .D(n36241), .Z(x_result_31__N_626[21])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32790_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32806_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[29]), 
         .D(n36265), .Z(x_result_31__N_626[29])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32806_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32796_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[24]), 
         .D(n36250), .Z(x_result_31__N_626[24])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32796_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32770_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[4]), 
         .D(n36190), .Z(x_result_31__N_626[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32770_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32782_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[17]), 
         .D(n36229), .Z(x_result_31__N_626[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32782_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32764_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[0]), 
         .D(n36175), .Z(x_result_31__N_626[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32764_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32788_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[20]), 
         .D(n36238), .Z(x_result_31__N_626[20])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32788_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32804_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[28]), 
         .D(n36262), .Z(x_result_31__N_626[28])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32804_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32798_3_lut_4_lut (.A(x_result_sel_add_x), .B(n41444), .C(x_result_31__N_1076[25]), 
         .D(n36253), .Z(x_result_31__N_626[25])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam i32798_3_lut_4_lut.init = 16'hf1e0;
    FD1P3DX store_operand_x_i0_i1 (.D(bypass_data_1[1]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i1.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i2 (.D(bypass_data_1[2]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i2.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i3 (.D(bypass_data_1[3]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i3.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i4 (.D(bypass_data_1[4]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i4.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i5 (.D(bypass_data_1[5]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i5.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i6 (.D(bypass_data_1[6]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i6.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i7 (.D(bypass_data_1[7]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i7.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i8 (.D(bypass_data_1[8]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[8])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i8.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i9 (.D(bypass_data_1[9]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[9])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i9.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i10 (.D(bypass_data_1[10]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[10])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i10.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i11 (.D(bypass_data_1[11]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[11])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i11.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i12 (.D(bypass_data_1[12]), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[12])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i12.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i13 (.D(bypass_data_1[13]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[13])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i13.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i14 (.D(bypass_data_1[14]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[14])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i14.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i15 (.D(bypass_data_1[15]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[15])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i15.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i16 (.D(bypass_data_1[16]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i16.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i17 (.D(bypass_data_1[17]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i17.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i18 (.D(bypass_data_1[18]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i18.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i19 (.D(bypass_data_1[19]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i19.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i20 (.D(bypass_data_1[20]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i20.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i21 (.D(bypass_data_1[21]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i21.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i22 (.D(bypass_data_1[22]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i22.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i23 (.D(bypass_data_1[23]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i23.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i24 (.D(bypass_data_1[24]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i24.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i25 (.D(bypass_data_1[25]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i25.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i26 (.D(bypass_data_1[26]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i26.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i27 (.D(bypass_data_1[27]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i27.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i28 (.D(bypass_data_1[28]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i28.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i29 (.D(bypass_data_1[29]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i29.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i30 (.D(bypass_data_1[30]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i30.GSR = "ENABLED";
    FD1P3DX store_operand_x_i0_i31 (.D(bypass_data_1[31]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_operand_x[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i31.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i3 (.D(branch_target_x_31__N_1120[1]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i3.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i4 (.D(branch_target_x_31__N_1120[2]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i4.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i5 (.D(branch_target_x_31__N_1120[3]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i5.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i6 (.D(branch_target_x_31__N_1120[4]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i6.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i7 (.D(branch_target_x_31__N_1120[5]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i7.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i8 (.D(branch_target_x_31__N_1120[6]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[8])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i8.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i9 (.D(branch_target_x_31__N_1120[7]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[9])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i9.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i10 (.D(branch_target_x_31__N_1120[8]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[10])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i10.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i11 (.D(branch_target_x_31__N_1120[9]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[11])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i11.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i12 (.D(branch_target_x_31__N_1120[10]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[12])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i12.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i13 (.D(branch_target_x_31__N_1120[11]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[13])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i13.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i14 (.D(branch_target_x_31__N_1120[12]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[14])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i14.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i15 (.D(branch_target_x_31__N_1120[13]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[15])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i15.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i16 (.D(branch_target_x_31__N_1120[14]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i16.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i17 (.D(branch_target_x_31__N_1120[15]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i17.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i18 (.D(branch_target_x_31__N_1120[16]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i18.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i19 (.D(branch_target_x_31__N_1120[17]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i19.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i20 (.D(branch_target_x_31__N_1120[18]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i20.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i21 (.D(branch_target_x_31__N_1120[19]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i21.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i22 (.D(branch_target_x_31__N_1120[20]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i22.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i23 (.D(branch_target_x_31__N_1120[21]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i23.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i24 (.D(branch_target_x_31__N_1120[22]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i24.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i25 (.D(branch_target_x_31__N_1120[23]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i25.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i26 (.D(branch_target_x_31__N_1120[24]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i26.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i27 (.D(branch_target_x_31__N_1120[25]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i27.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i28 (.D(branch_target_x_31__N_1120[26]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i28.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i29 (.D(branch_target_x_31__N_1120[27]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i29.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i30 (.D(branch_target_x_31__N_1120[28]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i30.GSR = "ENABLED";
    FD1P3DX branch_target_x_i2_i31 (.D(branch_target_x_31__N_1120[29]), .SP(REF_CLK_c_enable_823), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_x[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i31.GSR = "ENABLED";
    FD1P3DX csr_x_i0_i1 (.D(n41354), .SP(REF_CLK_c_enable_823), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(csr_x[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam csr_x_i0_i1.GSR = "ENABLED";
    FD1P3DX csr_x_i0_i2 (.D(n41351), .SP(REF_CLK_c_enable_823), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(csr_x[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam csr_x_i0_i2.GSR = "ENABLED";
    FD1P3DX csr_x_i0_i3 (.D(n41353), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(csr_x[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam csr_x_i0_i3.GSR = "ENABLED";
    FD1P3DX csr_x_i0_i4 (.D(n41352), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(csr_x[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam csr_x_i0_i4.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i3 (.D(branch_target_m_31__N_1167[1]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i3.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i4 (.D(branch_target_m_31__N_1167[2]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i4.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i5 (.D(branch_target_m_31__N_1167[3]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i5.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i6 (.D(branch_target_m_31__N_1167[4]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i6.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i7 (.D(branch_target_m_31__N_1167[5]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i7.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i8 (.D(branch_target_m_31__N_1167[6]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[8])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i8.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i9 (.D(branch_target_m_31__N_1167[7]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[9])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i9.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i10 (.D(branch_target_m_31__N_1167[8]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[10])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i10.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i11 (.D(branch_target_m_31__N_1167[9]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[11])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i11.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i12 (.D(branch_target_m_31__N_1167[10]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[12])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i12.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i13 (.D(branch_target_m_31__N_1167[11]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[13])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i13.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i14 (.D(branch_target_m_31__N_1167[12]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[14])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i14.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i15 (.D(branch_target_m_31__N_1167[13]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[15])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i15.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i16 (.D(branch_target_m_31__N_1167[14]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i16.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i17 (.D(branch_target_m_31__N_1167[15]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i17.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i18 (.D(branch_target_m_31__N_1167[16]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i18.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i19 (.D(branch_target_m_31__N_1167[17]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i19.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i20 (.D(branch_target_m_31__N_1167[18]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i20.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i21 (.D(branch_target_m_31__N_1167[19]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i21.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i22 (.D(branch_target_m_31__N_1167[20]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i22.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i23 (.D(branch_target_m_31__N_1167[21]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i23.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i24 (.D(branch_target_m_31__N_1167[22]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i24.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i25 (.D(branch_target_m_31__N_1167[23]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i25.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i26 (.D(branch_target_m_31__N_1167[24]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i26.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i27 (.D(branch_target_m_31__N_1167[25]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i27.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i28 (.D(branch_target_m_31__N_1167[26]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i28.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i29 (.D(branch_target_m_31__N_1167[27]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i29.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i30 (.D(branch_target_m_31__N_1167[28]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i30.GSR = "ENABLED";
    FD1P3DX branch_target_m_i2_i31 (.D(branch_target_m_31__N_1167[29]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(branch_target_m[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i31.GSR = "ENABLED";
    FD1P3DX eba_i8_i9 (.D(operand_1_x[9]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[9])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i9.GSR = "ENABLED";
    FD1P3DX eba_i8_i10 (.D(operand_1_x[10]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[10])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i10.GSR = "ENABLED";
    FD1P3DX eba_i8_i11 (.D(operand_1_x[11]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[11])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i11.GSR = "ENABLED";
    FD1P3DX eba_i8_i12 (.D(operand_1_x[12]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[12])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i12.GSR = "ENABLED";
    FD1P3DX eba_i8_i13 (.D(operand_1_x[13]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[13])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i13.GSR = "ENABLED";
    FD1P3DX eba_i8_i14 (.D(operand_1_x[14]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[14])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i14.GSR = "ENABLED";
    FD1P3BX eba_i8_i15 (.D(operand_1_x[15]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(eba[15])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i15.GSR = "ENABLED";
    FD1P3DX eba_i8_i16 (.D(operand_1_x[16]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i16.GSR = "ENABLED";
    FD1P3DX eba_i8_i17 (.D(operand_1_x[17]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i17.GSR = "ENABLED";
    FD1P3DX eba_i8_i18 (.D(operand_1_x[18]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i18.GSR = "ENABLED";
    FD1P3DX eba_i8_i19 (.D(operand_1_x[19]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i19.GSR = "ENABLED";
    FD1P3DX eba_i8_i20 (.D(operand_1_x[20]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i20.GSR = "ENABLED";
    FD1P3DX eba_i8_i21 (.D(operand_1_x[21]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i21.GSR = "ENABLED";
    FD1P3DX eba_i8_i22 (.D(operand_1_x[22]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i22.GSR = "ENABLED";
    FD1P3DX eba_i8_i23 (.D(operand_1_x[23]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i23.GSR = "ENABLED";
    FD1P3DX eba_i8_i24 (.D(operand_1_x[24]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i24.GSR = "ENABLED";
    FD1P3DX eba_i8_i25 (.D(operand_1_x[25]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i25.GSR = "ENABLED";
    FD1P3DX eba_i8_i26 (.D(operand_1_x[26]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i26.GSR = "ENABLED";
    FD1P3DX eba_i8_i27 (.D(operand_1_x[27]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i27.GSR = "ENABLED";
    FD1P3DX eba_i8_i28 (.D(operand_1_x[28]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i28.GSR = "ENABLED";
    FD1P3DX eba_i8_i29 (.D(operand_1_x[29]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i29.GSR = "ENABLED";
    FD1P3DX eba_i8_i30 (.D(operand_1_x[30]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i30.GSR = "ENABLED";
    FD1P3DX eba_i8_i31 (.D(operand_1_x[31]), .SP(eba_31__N_1111), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eba[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i31.GSR = "ENABLED";
    FD1S3DX operand_w_i1 (.D(operand_w_31__N_850[1]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(operand_w[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i1.GSR = "ENABLED";
    FD1S3DX operand_w_i2 (.D(operand_w_31__N_850[2]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(operand_w[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i2.GSR = "ENABLED";
    FD1S3DX operand_w_i3 (.D(operand_w_31__N_850[3]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(operand_w[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i3.GSR = "ENABLED";
    FD1S3DX operand_w_i4 (.D(operand_w_31__N_850[4]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(operand_w[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i4.GSR = "ENABLED";
    FD1S3DX operand_w_i5 (.D(operand_w_31__N_850[5]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(operand_w[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i5.GSR = "ENABLED";
    FD1S3DX operand_w_i6 (.D(operand_w_31__N_850[6]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(operand_w[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i6.GSR = "ENABLED";
    FD1S3DX operand_w_i7 (.D(operand_w_31__N_850[7]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(operand_w[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i7.GSR = "ENABLED";
    FD1S3DX operand_w_i8 (.D(operand_w_31__N_850[8]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(operand_w[8])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i8.GSR = "ENABLED";
    FD1S3DX operand_w_i9 (.D(operand_w_31__N_850[9]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(operand_w[9])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i9.GSR = "ENABLED";
    FD1S3DX operand_w_i10 (.D(operand_w_31__N_850[10]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[10])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i10.GSR = "ENABLED";
    FD1S3DX operand_w_i11 (.D(operand_w_31__N_850[11]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[11])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i11.GSR = "ENABLED";
    FD1S3DX operand_w_i12 (.D(operand_w_31__N_850[12]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[12])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i12.GSR = "ENABLED";
    FD1S3DX operand_w_i13 (.D(operand_w_31__N_850[13]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[13])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i13.GSR = "ENABLED";
    FD1S3DX operand_w_i14 (.D(operand_w_31__N_850[14]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[14])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i14.GSR = "ENABLED";
    FD1S3DX operand_w_i15 (.D(operand_w_31__N_850[15]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[15])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i15.GSR = "ENABLED";
    FD1S3DX operand_w_i16 (.D(operand_w_31__N_850[16]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i16.GSR = "ENABLED";
    FD1S3DX operand_w_i17 (.D(operand_w_31__N_850[17]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i17.GSR = "ENABLED";
    FD1S3DX operand_w_i18 (.D(operand_w_31__N_850[18]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i18.GSR = "ENABLED";
    FD1S3DX operand_w_i19 (.D(operand_w_31__N_850[19]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i19.GSR = "ENABLED";
    FD1S3DX operand_w_i20 (.D(operand_w_31__N_850[20]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i20.GSR = "ENABLED";
    FD1S3DX operand_w_i21 (.D(operand_w_31__N_850[21]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i21.GSR = "ENABLED";
    FD1S3DX operand_w_i22 (.D(operand_w_31__N_850[22]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i22.GSR = "ENABLED";
    FD1S3DX operand_w_i23 (.D(operand_w_31__N_850[23]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i23.GSR = "ENABLED";
    FD1S3DX operand_w_i24 (.D(operand_w_31__N_850[24]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i24.GSR = "ENABLED";
    FD1S3DX operand_w_i25 (.D(operand_w_31__N_850[25]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i25.GSR = "ENABLED";
    FD1S3DX operand_w_i26 (.D(operand_w_31__N_850[26]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i26.GSR = "ENABLED";
    FD1S3DX operand_w_i27 (.D(operand_w_31__N_850[27]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i27.GSR = "ENABLED";
    FD1S3DX operand_w_i28 (.D(operand_w_31__N_850[28]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i28.GSR = "ENABLED";
    FD1S3DX operand_w_i29 (.D(operand_w_31__N_850[29]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i29.GSR = "ENABLED";
    FD1S3DX operand_w_i30 (.D(operand_w_31__N_850[30]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i30.GSR = "ENABLED";
    FD1S3DX operand_w_i31 (.D(operand_w_31__N_850[31]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(operand_w[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i31.GSR = "ENABLED";
    FD1S3DX write_idx_w_i1 (.D(write_idx_m[1]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(write_idx_w[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_w_i1.GSR = "ENABLED";
    FD1S3DX write_idx_w_i2 (.D(write_idx_m[2]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(write_idx_w[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_w_i2.GSR = "ENABLED";
    FD1S3DX write_idx_w_i3 (.D(write_idx_m[3]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(write_idx_w[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_w_i3.GSR = "ENABLED";
    FD1S3DX write_idx_w_i4 (.D(write_idx_m[4]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(write_idx_w[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_w_i4.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i3 (.D(pc_m[3]), .SP(memop_pc_w_31__N_1229), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i3.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i4 (.D(pc_m[4]), .SP(memop_pc_w_31__N_1229), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i4.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i5 (.D(pc_m[5]), .SP(memop_pc_w_31__N_1229), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i5.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i6 (.D(pc_m[6]), .SP(memop_pc_w_31__N_1229), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i6.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i7 (.D(pc_m[7]), .SP(memop_pc_w_31__N_1229), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i7.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i8 (.D(pc_m[8]), .SP(memop_pc_w_31__N_1229), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[8])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i8.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i9 (.D(pc_m[9]), .SP(memop_pc_w_31__N_1229), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[9])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i9.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i10 (.D(pc_m[10]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[10])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i10.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i11 (.D(pc_m[11]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[11])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i11.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i12 (.D(pc_m[12]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[12])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i12.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i13 (.D(pc_m[13]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[13])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i13.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i14 (.D(pc_m[14]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[14])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i14.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i15 (.D(pc_m[15]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[15])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i15.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i16 (.D(pc_m[16]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i16.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i17 (.D(pc_m[17]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i17.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i18 (.D(pc_m[18]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i18.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i19 (.D(pc_m[19]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i19.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i20 (.D(pc_m[20]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i20.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i21 (.D(pc_m[21]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i21.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i22 (.D(pc_m[22]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i22.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i23 (.D(pc_m[23]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i23.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i24 (.D(pc_m[24]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i24.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i25 (.D(pc_m[25]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i25.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i26 (.D(pc_m[26]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i26.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i27 (.D(pc_m[27]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i27.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i28 (.D(pc_m[28]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i28.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i29 (.D(pc_m[29]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i29.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i30 (.D(pc_m[30]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i30.GSR = "ENABLED";
    FD1P3DX memop_pc_w_i2_i31 (.D(pc_m[31]), .SP(memop_pc_w_31__N_1229), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(memop_pc_w[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i31.GSR = "ENABLED";
    FD1P3DX write_idx_m_i0_i1 (.D(write_idx_m_4__N_1162[1]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(write_idx_m[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_m_i0_i1.GSR = "ENABLED";
    FD1P3DX write_idx_m_i0_i2 (.D(write_idx_m_4__N_1162[2]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(write_idx_m[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_m_i0_i2.GSR = "ENABLED";
    FD1P3DX write_idx_m_i0_i3 (.D(write_idx_m_4__N_1162[3]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(write_idx_m[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_m_i0_i3.GSR = "ENABLED";
    FD1P3DX write_idx_m_i0_i4 (.D(write_idx_m_4__N_1162[4]), .SP(REF_CLK_c_enable_1050), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(write_idx_m[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_m_i0_i4.GSR = "ENABLED";
    PFUMX i12658 (.BLUT(n17970), .ALUT(n17971), .C0(n37174), .Z(n17972));
    LUT4 operand_w_31__I_0_i5_3_lut (.A(operand_w[4]), .B(multiplier_result_w[4]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i6_3_lut (.A(operand_w[5]), .B(multiplier_result_w[5]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i7_3_lut (.A(operand_w[6]), .B(multiplier_result_w[6]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i8_3_lut (.A(operand_w[7]), .B(multiplier_result_w[7]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i17_3_lut (.A(operand_w[16]), .B(multiplier_result_w[16]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i17_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i18_3_lut (.A(operand_w[17]), .B(multiplier_result_w[17]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i18_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i19_3_lut (.A(operand_w[18]), .B(multiplier_result_w[18]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i19_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i20_3_lut (.A(operand_w[19]), .B(multiplier_result_w[19]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i20_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i21_3_lut (.A(operand_w[20]), .B(multiplier_result_w[20]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i21_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i22_3_lut (.A(operand_w[21]), .B(multiplier_result_w[21]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i22_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i23_3_lut (.A(operand_w[22]), .B(multiplier_result_w[22]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i23_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i24_3_lut (.A(operand_w[23]), .B(multiplier_result_w[23]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i24_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i25_3_lut (.A(operand_w[24]), .B(multiplier_result_w[24]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i25_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i26_3_lut (.A(operand_w[25]), .B(multiplier_result_w[25]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i26_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i27_3_lut (.A(operand_w[26]), .B(multiplier_result_w[26]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i27_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i28_3_lut (.A(operand_w[27]), .B(multiplier_result_w[27]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i28_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i29_3_lut (.A(operand_w[28]), .B(multiplier_result_w[28]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i29_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i30_3_lut (.A(operand_w[29]), .B(multiplier_result_w[29]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i30_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i31_3_lut (.A(operand_w[30]), .B(multiplier_result_w[30]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i31_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i32_3_lut (.A(operand_w[31]), .B(multiplier_result_w[31]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i32_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_1134 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_446)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1134.init = 16'h0f0e;
    LUT4 i15371_4_lut (.A(bie), .B(n31825), .C(im[2]), .D(csr_x[0]), 
         .Z(n5814[2])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15371_4_lut.init = 16'hc088;
    LUT4 i4387_4_lut (.A(im[8]), .B(deba[8]), .C(n41391), .D(n41288), 
         .Z(n5814[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4387_4_lut.init = 16'hcac0;
    FD1P3DX x_result_sel_sext_x_673 (.D(n31494), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(x_result_sel_sext_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam x_result_sel_sext_x_673.GSR = "ENABLED";
    FD1P3DX x_result_sel_mc_arith_x_672 (.D(n12412), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(x_result_sel_mc_arith_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam x_result_sel_mc_arith_x_672.GSR = "ENABLED";
    FD1P3DX w_result_sel_load_m_708 (.D(n12410), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(w_result_sel_load_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam w_result_sel_load_m_708.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_603 (.A(branch_flushX_m_N_1312), .B(n7_adj_6195), 
         .C(n30493), .D(n41420), .Z(branch_flushX_m)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_603.init = 16'h0200;
    FD1P3DX exception_m_714 (.D(n31804), .SP(REF_CLK_c_enable_1235), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(exception_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam exception_m_714.GSR = "ENABLED";
    LUT4 branch_flushX_m_I_49_4_lut (.A(condition_met_m), .B(exception_m), 
         .C(n30085), .D(n41450), .Z(branch_flushX_m_N_1312)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1677[29] 1687[9])
    defparam branch_flushX_m_I_49_4_lut.init = 16'hfcec;
    LUT4 i1_2_lut_adj_604 (.A(valid_m), .B(branch_m), .Z(n30085)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1677[37] 1678[55])
    defparam i1_2_lut_adj_604.init = 16'h8888;
    LUT4 i4401_4_lut (.A(im[15]), .B(deba[15]), .C(n41391), .D(n41288), 
         .Z(n5814[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4401_4_lut.init = 16'hcac0;
    LUT4 i4403_4_lut (.A(im[16]), .B(deba[16]), .C(n41391), .D(n41288), 
         .Z(n5814[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4403_4_lut.init = 16'hcac0;
    LUT4 i4405_4_lut (.A(im[17]), .B(deba[17]), .C(n41391), .D(n41288), 
         .Z(n5814[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4405_4_lut.init = 16'hcac0;
    LUT4 i4407_4_lut (.A(im[18]), .B(deba[18]), .C(n41391), .D(n41288), 
         .Z(n5814[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4407_4_lut.init = 16'hcac0;
    LUT4 n4_bdd_4_lut_4_lut (.A(operand_w[1]), .B(size_w[0]), .C(data_w[24]), 
         .D(data_w[8]), .Z(n41164)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam n4_bdd_4_lut_4_lut.init = 16'hfb40;
    LUT4 i4409_4_lut (.A(im[19]), .B(deba[19]), .C(n41391), .D(n41288), 
         .Z(n5814[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4409_4_lut.init = 16'hcac0;
    LUT4 n4_bdd_4_lut_34350_4_lut (.A(operand_w[1]), .B(size_w[0]), .C(data_w[25]), 
         .D(data_w[9]), .Z(n41160)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam n4_bdd_4_lut_34350_4_lut.init = 16'hfb40;
    LUT4 i4411_4_lut (.A(im[20]), .B(deba[20]), .C(n41391), .D(n41288), 
         .Z(n5814[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4411_4_lut.init = 16'hcac0;
    LUT4 n4_bdd_4_lut_34345_4_lut (.A(operand_w[1]), .B(size_w[0]), .C(data_w[26]), 
         .D(data_w[10]), .Z(n41156)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam n4_bdd_4_lut_34345_4_lut.init = 16'hfb40;
    LUT4 i4413_4_lut (.A(im[21]), .B(deba[21]), .C(n41391), .D(n41288), 
         .Z(n5814[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4413_4_lut.init = 16'hcac0;
    LUT4 n4_bdd_4_lut_34340_4_lut (.A(operand_w[1]), .B(size_w[0]), .C(data_w[27]), 
         .D(data_w[11]), .Z(n41152)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam n4_bdd_4_lut_34340_4_lut.init = 16'hfb40;
    LUT4 i4415_4_lut (.A(im[22]), .B(deba[22]), .C(n41391), .D(n41288), 
         .Z(n5814[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4415_4_lut.init = 16'hcac0;
    LUT4 n4_bdd_4_lut_34335_4_lut (.A(operand_w[1]), .B(size_w[0]), .C(data_w[28]), 
         .D(data_w[12]), .Z(n41148)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam n4_bdd_4_lut_34335_4_lut.init = 16'hfb40;
    LUT4 i4417_4_lut (.A(im[23]), .B(deba[23]), .C(n41391), .D(n41288), 
         .Z(n5814[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4417_4_lut.init = 16'hcac0;
    LUT4 n4_bdd_4_lut_34330_4_lut (.A(operand_w[1]), .B(size_w[0]), .C(data_w[29]), 
         .D(data_w[13]), .Z(n41144)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam n4_bdd_4_lut_34330_4_lut.init = 16'hfb40;
    LUT4 operand_w_31__I_0_i2_3_lut (.A(operand_w[1]), .B(multiplier_result_w[1]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 i4419_4_lut (.A(im[24]), .B(deba[24]), .C(n41391), .D(n41288), 
         .Z(n5814[24])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4419_4_lut.init = 16'hcac0;
    LUT4 n4_bdd_4_lut_34325_4_lut (.A(operand_w[1]), .B(size_w[0]), .C(data_w[30]), 
         .D(data_w[14]), .Z(n41140)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam n4_bdd_4_lut_34325_4_lut.init = 16'hfb40;
    LUT4 i4421_4_lut (.A(im[25]), .B(deba[25]), .C(n41391), .D(n41288), 
         .Z(n5814[25])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4421_4_lut.init = 16'hcac0;
    LUT4 n4_bdd_4_lut_34320_4_lut (.A(operand_w[1]), .B(size_w[0]), .C(data_w[31]), 
         .D(data_w[15]), .Z(n41136)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam n4_bdd_4_lut_34320_4_lut.init = 16'hfb40;
    LUT4 i4423_4_lut (.A(im[26]), .B(deba[26]), .C(n41391), .D(n41288), 
         .Z(n5814[26])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4423_4_lut.init = 16'hcac0;
    LUT4 n41730_bdd_3_lut (.A(n41730), .B(n41728), .C(x_result_sel_sext_x), 
         .Z(n41731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41730_bdd_3_lut.init = 16'hcaca;
    LUT4 i4425_4_lut (.A(im[27]), .B(deba[27]), .C(n41391), .D(n41288), 
         .Z(n5814[27])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4425_4_lut.init = 16'hcac0;
    LUT4 i4427_4_lut (.A(im[28]), .B(deba[28]), .C(n41391), .D(n41288), 
         .Z(n5814[28])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4427_4_lut.init = 16'hcac0;
    LUT4 mux_508_i29_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[30]), .C(eba[30]), 
         .Z(n41502)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i29_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 i4429_4_lut (.A(im[29]), .B(deba[29]), .C(n41391), .D(n41288), 
         .Z(n5814[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4429_4_lut.init = 16'hcac0;
    LUT4 mux_508_i29_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[30]), .C(branch_target_x[30]), 
         .Z(n41501)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i29_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 i4431_4_lut (.A(im[30]), .B(deba[30]), .C(n41391), .D(n41288), 
         .Z(n5814[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4431_4_lut.init = 16'hcac0;
    LUT4 logic_result_x_8__bdd_4_lut_34551 (.A(size_x[1]), .B(size_x[0]), 
         .C(operand_0_x[8]), .D(operand_0_x[7]), .Z(n41728)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam logic_result_x_8__bdd_4_lut_34551.init = 16'hf1e0;
    LUT4 i4433_4_lut (.A(im[31]), .B(deba[31]), .C(n41391), .D(n41288), 
         .Z(n5814[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i4433_4_lut.init = 16'hcac0;
    LUT4 mux_508_i28_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[29]), .C(eba[29]), 
         .Z(n41505)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i28_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i28_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[29]), .C(branch_target_x[29]), 
         .Z(n41504)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i28_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 i1_2_lut_rep_1135 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_445)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1135.init = 16'h0f0e;
    LUT4 mux_508_i27_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[28]), .C(eba[28]), 
         .Z(n41508)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i27_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i27_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[28]), .C(branch_target_x[28]), 
         .Z(n41507)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i27_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 i1_2_lut_rep_1136 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_444)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1136.init = 16'h0f0e;
    LUT4 mux_508_i26_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[27]), .C(eba[27]), 
         .Z(n41511)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i26_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i26_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[27]), .C(branch_target_x[27]), 
         .Z(n41510)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i26_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 logic_result_x_8__bdd_4_lut_34502 (.A(n5814[8]), .B(n41168), .C(n5915), 
         .D(csr_x[2]), .Z(n41727)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C (D)))) */ ;
    defparam logic_result_x_8__bdd_4_lut_34502.init = 16'hc0a0;
    LUT4 mux_508_i25_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[26]), .C(eba[26]), 
         .Z(n41514)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i25_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 i1_3_lut_4_lut_adj_605 (.A(n45175), .B(REF_CLK_c_enable_388), .C(n35639), 
         .D(n31334), .Z(n31279)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_605.init = 16'h0008;
    LUT4 mux_508_i25_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[26]), .C(branch_target_x[26]), 
         .Z(n41513)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i25_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i24_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[25]), .C(eba[25]), 
         .Z(n41517)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i24_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i24_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[25]), .C(branch_target_x[25]), 
         .Z(n41516)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i24_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 i1_3_lut_rep_1137 (.A(state[2]), .B(state_adj_6256[1]), .C(n30493), 
         .D(n7_adj_6195), .Z(n45171)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_rep_1137.init = 16'h0008;
    LUT4 mux_508_i23_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[24]), .C(eba[24]), 
         .Z(n41520)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i23_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i23_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[24]), .C(branch_target_x[24]), 
         .Z(n41519)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i23_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 i1_3_lut_rep_1138 (.A(state[2]), .B(state_adj_6256[1]), .C(n30493), 
         .D(n7_adj_6195), .Z(REF_CLK_c_enable_1235)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_rep_1138.init = 16'h0008;
    LUT4 mux_508_i22_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[23]), .C(eba[23]), 
         .Z(n41523)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i22_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i22_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[23]), .C(branch_target_x[23]), 
         .Z(n41522)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i22_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 i1_3_lut_rep_1139 (.A(state[2]), .B(state_adj_6256[1]), .C(n30493), 
         .D(n7_adj_6195), .Z(REF_CLK_c_enable_1050)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_rep_1139.init = 16'h0008;
    LUT4 mux_508_i21_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[22]), .C(eba[22]), 
         .Z(n41526)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i21_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i21_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[22]), .C(branch_target_x[22]), 
         .Z(n41525)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i21_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i20_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[21]), .C(eba[21]), 
         .Z(n41529)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i20_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i20_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[21]), .C(branch_target_x[21]), 
         .Z(n41528)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i20_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 n41737_bdd_3_lut (.A(n41737), .B(n41735), .C(x_result_sel_sext_x), 
         .Z(n41738)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41737_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_508_i19_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[20]), .C(eba[20]), 
         .Z(n41532)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i19_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i19_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[20]), .C(branch_target_x[20]), 
         .Z(n41531)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i19_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 i1_3_lut_rep_1140 (.A(state[2]), .B(state_adj_6256[1]), .C(n30493), 
         .D(n7_adj_6195), .Z(REF_CLK_c_enable_1299)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_rep_1140.init = 16'h0008;
    LUT4 mux_508_i18_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[19]), .C(eba[19]), 
         .Z(n41535)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i18_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i18_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[19]), .C(branch_target_x[19]), 
         .Z(n41534)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i18_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i17_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[18]), .C(eba[18]), 
         .Z(n41538)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i17_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i17_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[18]), .C(branch_target_x[18]), 
         .Z(n41537)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i17_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 n41739_bdd_3_lut (.A(n41739), .B(adder_result_x[9]), .C(x_result_sel_add_x), 
         .Z(x_result[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41739_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_508_i16_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[17]), .C(eba[17]), 
         .Z(n41541)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i16_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i16_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[17]), .C(branch_target_x[17]), 
         .Z(n41540)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i16_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 logic_result_x_10__bdd_4_lut_34512 (.A(n39321), .B(n5915), .C(n39320), 
         .D(csr_x[2]), .Z(n41741)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam logic_result_x_10__bdd_4_lut_34512.init = 16'hc088;
    LUT4 mux_508_i15_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[16]), .C(eba[16]), 
         .Z(n41544)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i15_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 i1_3_lut_4_lut_adj_606 (.A(n41205), .B(n30070), .C(n15), .D(n41197), 
         .Z(stall_a)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1873[20] 1904[21])
    defparam i1_3_lut_4_lut_adj_606.init = 16'hfff8;
    LUT4 mux_508_i15_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[16]), .C(branch_target_x[16]), 
         .Z(n41543)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i15_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 logic_result_x_10__bdd_4_lut_35767 (.A(size_x[1]), .B(size_x[0]), 
         .C(operand_0_x[10]), .D(operand_0_x[7]), .Z(n41742)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam logic_result_x_10__bdd_4_lut_35767.init = 16'hf1e0;
    LUT4 mux_3055_i7_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra [6]), 
         .D(adder_result_x[8]), .Z(n7388[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3055_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_4_lut_adj_607 (.A(n41232), .B(REF_CLK_c_enable_388), .C(n41233), 
         .D(n34890), .Z(deba_31__N_1118)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_607.init = 16'h0800;
    LUT4 mux_508_i14_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[15]), .C(eba[15]), 
         .Z(n41547)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i14_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i14_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[15]), .C(branch_target_x[15]), 
         .Z(n41546)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i14_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 logic_result_x_10__bdd_3_lut_35768 (.A(size_x[1]), .B(size_x[0]), 
         .C(operand_0_x[10]), .Z(n41743)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam logic_result_x_10__bdd_3_lut_35768.init = 16'hacac;
    LUT4 i1_2_lut_rep_1096 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_434)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1096.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_1097 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_433)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1097.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_1098 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_432)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1098.init = 16'h0f0e;
    LUT4 mux_76_i1_3_lut (.A(n1261[0]), .B(adder_result_x[0]), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i1_3_lut.init = 16'hcaca;
    LUT4 mux_508_i13_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[14]), .C(eba[14]), 
         .Z(n41550)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i13_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i13_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[14]), .C(branch_target_x[14]), 
         .Z(n41549)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i13_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 mux_76_i2_3_lut (.A(n1261[1]), .B(adder_result_x[1]), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_1141 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(n45175)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1141.init = 16'h0f0e;
    LUT4 mux_76_i3_3_lut (.A(n1261[2]), .B(adder_result_x[2]), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i3_3_lut.init = 16'hcaca;
    LUT4 mux_76_i5_3_lut (.A(n1261[4]), .B(adder_result_x[4]), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i5_3_lut.init = 16'hcaca;
    LUT4 mux_508_i12_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[13]), .C(eba[13]), 
         .Z(n41553)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i12_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_76_i6_3_lut (.A(n1261[5]), .B(adder_result_x[5]), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i6_3_lut.init = 16'hcaca;
    LUT4 mux_508_i12_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[13]), .C(branch_target_x[13]), 
         .Z(n41552)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i12_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 mux_76_i7_3_lut (.A(n1261[6]), .B(adder_result_x[6]), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i7_3_lut.init = 16'hcaca;
    LUT4 mux_76_i8_3_lut (.A(n1261[7]), .B(adder_result_x[7]), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i8_3_lut.init = 16'hcaca;
    LUT4 mux_2953_i2_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7206), .D(adder_result_x[3]), 
         .Z(n7190[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2953_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 n10760_bdd_4_lut_33731 (.A(n41288), .B(n41391), .C(im[13]), .D(deba[13]), 
         .Z(n39330)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (D))) */ ;
    defparam n10760_bdd_4_lut_33731.init = 16'hec20;
    LUT4 mux_76_i16_3_lut (.A(n1261[15]), .B(adder_result_x[15]), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i16_3_lut.init = 16'hcaca;
    LUT4 mux_508_i11_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[12]), .C(eba[12]), 
         .Z(n41556)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i11_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_76_i17_3_lut (.A(n1261[16]), .B(\adder_result_x[16] ), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i17_3_lut.init = 16'hcaca;
    LUT4 mux_508_i11_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[12]), .C(branch_target_x[12]), 
         .Z(n41555)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i11_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 mux_76_i18_3_lut (.A(n1261[17]), .B(\adder_result_x[17] ), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i18_3_lut.init = 16'hcaca;
    LUT4 n41744_bdd_3_lut (.A(n41744), .B(n41742), .C(x_result_sel_sext_x), 
         .Z(n41745)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41744_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_76_i19_3_lut (.A(n1261[18]), .B(\adder_result_x[18] ), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i19_3_lut.init = 16'hcaca;
    LUT4 mux_508_i10_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[11]), .C(eba[11]), 
         .Z(n41559)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i10_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_76_i20_3_lut (.A(n1261[19]), .B(\adder_result_x[19] ), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i20_3_lut.init = 16'hcaca;
    LUT4 mux_508_i10_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[11]), .C(branch_target_x[11]), 
         .Z(n41558)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i10_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 mux_76_i21_3_lut (.A(n1261[20]), .B(\adder_result_x[20] ), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i21_3_lut.init = 16'hcaca;
    LUT4 mux_3021_i5_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7344), .D(adder_result_x[6]), 
         .Z(n7322[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3021_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_rep_1142 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_1624)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1142.init = 16'h0f0e;
    LUT4 mux_76_i22_3_lut (.A(n1261[21]), .B(\adder_result_x[21] ), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i22_3_lut.init = 16'hcaca;
    LUT4 mux_76_i23_3_lut (.A(n1261[22]), .B(\adder_result_x[22] ), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i23_3_lut.init = 16'hcaca;
    LUT4 mux_508_i9_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[10]), .C(eba[10]), 
         .Z(n41562)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i9_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_76_i24_3_lut (.A(n1261[23]), .B(\adder_result_x[23] ), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i24_3_lut.init = 16'hcaca;
    LUT4 mux_508_i9_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[10]), .C(branch_target_x[10]), 
         .Z(n41561)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i9_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 mux_76_i25_3_lut (.A(n1261[24]), .B(\adder_result_x[24] ), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i25_3_lut.init = 16'hcaca;
    LUT4 mux_76_i26_3_lut (.A(n1261[25]), .B(\adder_result_x[25] ), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i26_3_lut.init = 16'hcaca;
    LUT4 mux_76_i27_3_lut (.A(n1261[26]), .B(\adder_result_x[26] ), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i27_3_lut.init = 16'hcaca;
    LUT4 mux_508_i8_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[9]), .C(eba[9]), 
         .Z(n41565)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i8_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_76_i28_3_lut (.A(n1261[27]), .B(\adder_result_x[27] ), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i28_3_lut.init = 16'hcaca;
    LUT4 mux_508_i8_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[9]), .C(branch_target_x[9]), 
         .Z(n41564)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i8_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 mux_76_i29_3_lut (.A(n1261[28]), .B(\adder_result_x[28] ), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i29_3_lut.init = 16'hcaca;
    LUT4 n41746_bdd_3_lut (.A(n41746), .B(adder_result_x[10]), .C(x_result_sel_add_x), 
         .Z(x_result[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41746_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_76_i30_3_lut (.A(n1261[29]), .B(\adder_result_x[29] ), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i30_3_lut.init = 16'hcaca;
    LUT4 mux_76_i31_3_lut (.A(n1261[30]), .B(\adder_result_x[30] ), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i31_3_lut.init = 16'hcaca;
    LUT4 mux_508_i7_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[8]), .C(eba[8]), 
         .Z(n41568)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i7_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_76_i32_3_lut (.A(n1261[31]), .B(\adder_result_x[31] ), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i32_3_lut.init = 16'hcaca;
    LUT4 mux_508_i7_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[8]), .C(branch_target_x[8]), 
         .Z(n41567)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i7_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 logic_result_x_11__bdd_4_lut_34517 (.A(n39324), .B(n5915), .C(n39323), 
         .D(csr_x[2]), .Z(n41748)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam logic_result_x_11__bdd_4_lut_34517.init = 16'hc088;
    LUT4 mux_2987_i4_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7276), .D(adder_result_x[5]), 
         .Z(n7256[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2987_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i34316_then_3_lut (.A(csr_x[0]), .B(jrx_csr_read_data[4]), .C(csr_x[2]), 
         .Z(n41571)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i34316_then_3_lut.init = 16'h8080;
    LUT4 mux_2987_i3_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7274), .D(adder_result_x[4]), 
         .Z(n7256[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2987_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_2987_i2_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7272), .D(adder_result_x[3]), 
         .Z(n7256[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2987_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_2987_i1_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7270), .D(adder_result_x[2]), 
         .Z(n7256[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2987_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_rep_1143 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_823)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1143.init = 16'h0f0e;
    LUT4 mux_2953_i9_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7220), .D(adder_result_x[10]), 
         .Z(n7190[8])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2953_i9_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i34316_else_3_lut (.A(csr_x[0]), .B(n41308), .C(im[4]), .D(csr_x[2]), 
         .Z(n41570)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i34316_else_3_lut.init = 16'h0020;
    LUT4 mux_3021_i11_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7356), 
         .D(adder_result_x[12]), .Z(n7322[10])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3021_i11_3_lut_4_lut.init = 16'hf4b0;
    LUT4 logic_result_x_11__bdd_4_lut_35539 (.A(size_x[1]), .B(size_x[0]), 
         .C(operand_0_x[11]), .D(operand_0_x[7]), .Z(n41749)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam logic_result_x_11__bdd_4_lut_35539.init = 16'hf1e0;
    LUT4 mux_3021_i10_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7354), 
         .D(adder_result_x[11]), .Z(n7322[9])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3021_i10_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3021_i9_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7352), .D(adder_result_x[10]), 
         .Z(n7322[8])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3021_i9_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_76_i4_3_lut (.A(n1261[3]), .B(adder_result_x[3]), .C(x_result_sel_add_x), 
         .Z(x_result_31__N_1076[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i4_3_lut.init = 16'hcaca;
    LUT4 i34312_then_3_lut (.A(csr_x[0]), .B(jrx_csr_read_data[5]), .C(csr_x[2]), 
         .Z(n41574)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i34312_then_3_lut.init = 16'h8080;
    LUT4 i34312_else_3_lut (.A(csr_x[0]), .B(n41308), .C(im[5]), .D(csr_x[2]), 
         .Z(n41573)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i34312_else_3_lut.init = 16'h0020;
    LUT4 logic_result_x_11__bdd_3_lut_35540 (.A(size_x[1]), .B(size_x[0]), 
         .C(operand_0_x[11]), .Z(n41750)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam logic_result_x_11__bdd_3_lut_35540.init = 16'hacac;
    LUT4 mux_3021_i8_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7350), .D(adder_result_x[9]), 
         .Z(n7322[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3021_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_rep_1144 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_1030)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1144.init = 16'h0f0e;
    LUT4 i1_3_lut_rep_1147 (.A(n41232), .B(n41233), .C(n15), .D(n41196), 
         .Z(n45181)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_3_lut_rep_1147.init = 16'h0002;
    LUT4 mux_3021_i7_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7348), .D(adder_result_x[8]), 
         .Z(n7322[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3021_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_3_lut_rep_1148 (.A(n41232), .B(n41233), .C(n15), .D(n41196), 
         .Z(REF_CLK_c_enable_1178)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_3_lut_rep_1148.init = 16'h0002;
    LUT4 mux_3021_i6_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7346), .D(adder_result_x[7]), 
         .Z(n7322[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3021_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3021_i4_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7342), .D(adder_result_x[5]), 
         .Z(n7322[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3021_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_3_lut_4_lut_rep_1149 (.A(n41205), .B(n30070), .C(n15), .D(n41197), 
         .Z(n45183)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1873[20] 1904[21])
    defparam i1_3_lut_4_lut_rep_1149.init = 16'hfff8;
    LUT4 n4_bdd_3_lut_34322 (.A(operand_w[15]), .B(multiplier_result_w[15]), 
         .C(w_result_sel_mul_w), .Z(n41138)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n4_bdd_3_lut_34322.init = 16'hcaca;
    LUT4 stall_m_N_1151_I_0_797_rep_18_2_lut_4_lut (.A(n7_adj_6195), .B(n41420), 
         .C(n30493), .D(branch_flushX_m_N_1312), .Z(n30479)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam stall_m_N_1151_I_0_797_rep_18_2_lut_4_lut.init = 16'h0400;
    LUT4 bypass_data_0_31__I_14_i9_3_lut (.A(m_result[8]), .B(x_result[8]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i9_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_812_4_lut (.A(n7_adj_6195), .B(n41420), .C(n30493), 
         .D(n41283), .Z(n41217)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_rep_812_4_lut.init = 16'h0400;
    LUT4 i7019_2_lut_4_lut (.A(n7_adj_6195), .B(n41420), .C(n30493), .D(dcache_refill_request), 
         .Z(REF_CLK_c_enable_1513)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;
    defparam i7019_2_lut_4_lut.init = 16'hff04;
    LUT4 mux_46_i9_4_lut (.A(n7609[8]), .B(w_result[8]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i9_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i10_3_lut (.A(m_result[9]), .B(x_result[9]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i10_3_lut.init = 16'hcaca;
    LUT4 mux_46_i10_4_lut (.A(n7609[9]), .B(w_result[9]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i10_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i11_3_lut (.A(m_result[10]), .B(x_result[10]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i11_3_lut.init = 16'hcaca;
    LUT4 mux_46_i11_4_lut (.A(n7609[10]), .B(w_result[10]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i11_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i12_3_lut (.A(m_result[11]), .B(x_result[11]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i12_3_lut.init = 16'hcaca;
    LUT4 mux_46_i12_4_lut (.A(n7609[11]), .B(w_result[11]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i12_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i13_3_lut (.A(m_result[12]), .B(x_result[12]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i13_3_lut.init = 16'hcaca;
    LUT4 mux_46_i13_4_lut (.A(n7609[12]), .B(w_result[12]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i13_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i14_3_lut (.A(m_result[13]), .B(x_result[13]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i14_3_lut.init = 16'hcaca;
    FD1P3DX valid_m_665 (.D(n31655), .SP(REF_CLK_c_enable_1513), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(valid_m)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2264[5] 2299[8])
    defparam valid_m_665.GSR = "ENABLED";
    LUT4 mux_46_i14_4_lut (.A(n7609[13]), .B(w_result[13]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i14_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i15_3_lut (.A(m_result[14]), .B(x_result[14]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i15_3_lut.init = 16'hcaca;
    LUT4 mux_46_i15_4_lut (.A(n7609[14]), .B(w_result[14]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i15_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i9_3_lut (.A(m_result[8]), .B(x_result[8]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i9_3_lut.init = 16'hcaca;
    LUT4 mux_52_i9_4_lut (.A(n7677[8]), .B(w_result[8]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i9_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i10_3_lut (.A(m_result[9]), .B(x_result[9]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i10_3_lut.init = 16'hcaca;
    LUT4 mux_52_i10_4_lut (.A(n7677[9]), .B(w_result[9]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i10_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i11_3_lut (.A(m_result[10]), .B(x_result[10]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i11_3_lut.init = 16'hcaca;
    LUT4 mux_52_i11_4_lut (.A(n7677[10]), .B(w_result[10]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i11_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i12_3_lut (.A(m_result[11]), .B(x_result[11]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i12_3_lut.init = 16'hcaca;
    LUT4 mux_52_i12_4_lut (.A(n7677[11]), .B(w_result[11]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i12_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i13_3_lut (.A(m_result[12]), .B(x_result[12]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i13_3_lut.init = 16'hcaca;
    LUT4 mux_52_i13_4_lut (.A(n7677[12]), .B(w_result[12]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i13_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i14_3_lut (.A(m_result[13]), .B(x_result[13]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i14_3_lut.init = 16'hcaca;
    LUT4 mux_52_i14_4_lut (.A(n7677[13]), .B(w_result[13]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i14_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i15_3_lut (.A(m_result[14]), .B(x_result[14]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i15_3_lut.init = 16'hcaca;
    LUT4 mux_52_i15_4_lut (.A(n7677[14]), .B(w_result[14]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i15_4_lut.init = 16'hcac0;
    LUT4 i12659_3_lut (.A(n17972), .B(x_result[0]), .C(raw_x_0), .Z(bypass_data_0_31__N_882[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(707[6:13])
    defparam i12659_3_lut.init = 16'hcaca;
    LUT4 i12655_4_lut (.A(n7609[0]), .B(w_result[0]), .C(raw_w_0), .D(n6518), 
         .Z(n17969)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(709[6:13])
    defparam i12655_4_lut.init = 16'hcac0;
    LUT4 i12661_3_lut (.A(n17972), .B(x_result[0]), .C(raw_x_1), .Z(bypass_data_1_31__N_914[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(708[6:13])
    defparam i12661_3_lut.init = 16'hcaca;
    LUT4 i12660_4_lut (.A(n7677[0]), .B(w_result[0]), .C(raw_w_1), .D(n6648), 
         .Z(n17974)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(710[6:13])
    defparam i12660_4_lut.init = 16'hcac0;
    LUT4 i14165_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7338), .D(adder_result_x[3]), 
         .Z(n7322[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam i14165_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_rep_1086 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_729)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1086.init = 16'h0f0e;
    LUT4 i2_4_lut (.A(bus_error_f_N_1884), .B(stall_wb_load), .C(branch_m), 
         .D(exception_m), .Z(n7_adj_6195)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;
    defparam i2_4_lut.init = 16'heeec;
    LUT4 n10760_bdd_4_lut_33745 (.A(n41288), .B(n41391), .C(im[14]), .D(deba[14]), 
         .Z(n39333)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (D))) */ ;
    defparam n10760_bdd_4_lut_33745.init = 16'hec20;
    LUT4 mux_3055_i1_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra [0]), 
         .D(adder_result_x[2]), .Z(n7388[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3055_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3055_i2_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra [1]), 
         .D(adder_result_x[3]), .Z(n7388[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3055_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3021_i3_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7340), .D(adder_result_x[4]), 
         .Z(n7322[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3021_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3021_i1_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7336), .D(adder_result_x[2]), 
         .Z(n7322[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3021_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_46_i2_4_lut (.A(n7609[1]), .B(w_result[1]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i2_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i3_3_lut (.A(m_result[2]), .B(x_result[2]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i3_3_lut.init = 16'hcaca;
    LUT4 mux_46_i3_4_lut (.A(n7609[2]), .B(w_result[2]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i3_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i4_3_lut (.A(m_result[3]), .B(x_result[3]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i4_3_lut.init = 16'hcaca;
    LUT4 mux_46_i4_4_lut (.A(n7609[3]), .B(w_result[3]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i4_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i5_3_lut (.A(m_result[4]), .B(x_result[4]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i5_3_lut.init = 16'hcaca;
    LUT4 mux_46_i5_4_lut (.A(n7609[4]), .B(w_result[4]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i5_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i6_3_lut (.A(m_result[5]), .B(x_result[5]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i6_3_lut.init = 16'hcaca;
    LUT4 mux_46_i6_4_lut (.A(n7609[5]), .B(w_result[5]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i6_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i7_3_lut (.A(m_result[6]), .B(x_result[6]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i7_3_lut.init = 16'hcaca;
    LUT4 mux_46_i7_4_lut (.A(n7609[6]), .B(w_result[6]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i7_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i8_3_lut (.A(m_result[7]), .B(x_result[7]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i8_3_lut.init = 16'hcaca;
    LUT4 mux_46_i8_4_lut (.A(n7609[7]), .B(w_result[7]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i8_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i16_3_lut (.A(m_result[15]), .B(x_result[15]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i16_3_lut.init = 16'hcaca;
    LUT4 mux_46_i16_4_lut (.A(n7609[15]), .B(w_result[15]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i16_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i17_3_lut (.A(m_result[16]), .B(x_result[16]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i17_3_lut.init = 16'hcaca;
    LUT4 mux_46_i17_4_lut (.A(n7609[16]), .B(w_result[16]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i17_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i18_3_lut (.A(m_result[17]), .B(x_result[17]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i18_3_lut.init = 16'hcaca;
    LUT4 mux_2953_i3_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7208), .D(adder_result_x[4]), 
         .Z(n7190[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2953_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_46_i18_4_lut (.A(n7609[17]), .B(w_result[17]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i18_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i19_3_lut (.A(m_result[18]), .B(x_result[18]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i19_3_lut.init = 16'hcaca;
    LUT4 mux_46_i19_4_lut (.A(n7609[18]), .B(w_result[18]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i19_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i20_3_lut (.A(m_result[19]), .B(x_result[19]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i20_3_lut.init = 16'hcaca;
    LUT4 mux_46_i20_4_lut (.A(n7609[19]), .B(w_result[19]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i20_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i21_3_lut (.A(m_result[20]), .B(x_result[20]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i21_3_lut.init = 16'hcaca;
    LUT4 mux_46_i21_4_lut (.A(n7609[20]), .B(w_result[20]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i21_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i22_3_lut (.A(m_result[21]), .B(x_result[21]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i22_3_lut.init = 16'hcaca;
    LUT4 mux_46_i22_4_lut (.A(n7609[21]), .B(w_result[21]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i22_4_lut.init = 16'hcac0;
    LUT4 mux_3055_i5_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra [4]), 
         .D(adder_result_x[6]), .Z(n7388[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3055_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 bypass_data_0_31__I_14_i23_3_lut (.A(m_result[22]), .B(x_result[22]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i23_3_lut.init = 16'hcaca;
    LUT4 mux_46_i23_4_lut (.A(n7609[22]), .B(w_result[22]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i23_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i24_3_lut (.A(m_result[23]), .B(x_result[23]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i24_3_lut.init = 16'hcaca;
    LUT4 mux_46_i24_4_lut (.A(n7609[23]), .B(w_result[23]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i24_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i25_3_lut (.A(m_result[24]), .B(x_result[24]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i25_3_lut.init = 16'hcaca;
    LUT4 mux_46_i25_4_lut (.A(n7609[24]), .B(w_result[24]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[24])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i25_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i26_3_lut (.A(m_result[25]), .B(x_result[25]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i26_3_lut.init = 16'hcaca;
    LUT4 mux_46_i26_4_lut (.A(n7609[25]), .B(w_result[25]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[25])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i26_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i27_3_lut (.A(m_result[26]), .B(x_result[26]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i27_3_lut.init = 16'hcaca;
    LUT4 mux_46_i27_4_lut (.A(n7609[26]), .B(w_result[26]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[26])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i27_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i28_3_lut (.A(m_result[27]), .B(x_result[27]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i28_3_lut.init = 16'hcaca;
    LUT4 mux_46_i28_4_lut (.A(n7609[27]), .B(w_result[27]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[27])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i28_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i29_3_lut (.A(m_result[28]), .B(x_result[28]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i29_3_lut.init = 16'hcaca;
    LUT4 mux_46_i29_4_lut (.A(n7609[28]), .B(w_result[28]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[28])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i29_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i30_3_lut (.A(m_result[29]), .B(x_result[29]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i30_3_lut.init = 16'hcaca;
    LUT4 mux_46_i30_4_lut (.A(n7609[29]), .B(w_result[29]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i30_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i31_3_lut (.A(m_result[30]), .B(x_result[30]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i31_3_lut.init = 16'hcaca;
    LUT4 mux_46_i31_4_lut (.A(n7609[30]), .B(w_result[30]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i31_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_14_i32_3_lut (.A(m_result[31]), .B(x_result[31]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_882[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_14_i32_3_lut.init = 16'hcaca;
    LUT4 mux_46_i32_4_lut (.A(n7609[31]), .B(w_result[31]), .C(raw_w_0), 
         .D(n6518), .Z(bypass_data_0_31__N_1012[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i32_4_lut.init = 16'hcac0;
    LUT4 mux_52_i2_4_lut (.A(n7677[1]), .B(w_result[1]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i2_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i3_3_lut (.A(m_result[2]), .B(x_result[2]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i3_3_lut.init = 16'hcaca;
    LUT4 mux_52_i3_4_lut (.A(n7677[2]), .B(w_result[2]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i3_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i4_3_lut (.A(m_result[3]), .B(x_result[3]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i4_3_lut.init = 16'hcaca;
    LUT4 mux_52_i4_4_lut (.A(n7677[3]), .B(w_result[3]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i4_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i5_3_lut (.A(m_result[4]), .B(x_result[4]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i5_3_lut.init = 16'hcaca;
    LUT4 mux_52_i5_4_lut (.A(n7677[4]), .B(w_result[4]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i5_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i6_3_lut (.A(m_result[5]), .B(x_result[5]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i6_3_lut.init = 16'hcaca;
    LUT4 mux_52_i6_4_lut (.A(n7677[5]), .B(w_result[5]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i6_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i7_3_lut (.A(m_result[6]), .B(x_result[6]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i7_3_lut.init = 16'hcaca;
    LUT4 mux_52_i7_4_lut (.A(n7677[6]), .B(w_result[6]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i7_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i8_3_lut (.A(m_result[7]), .B(x_result[7]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i8_3_lut.init = 16'hcaca;
    LUT4 mux_52_i8_4_lut (.A(n7677[7]), .B(w_result[7]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i8_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i16_3_lut (.A(m_result[15]), .B(x_result[15]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i16_3_lut.init = 16'hcaca;
    LUT4 mux_52_i16_4_lut (.A(n7677[15]), .B(w_result[15]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i16_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i17_3_lut (.A(m_result[16]), .B(x_result[16]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i17_3_lut.init = 16'hcaca;
    LUT4 mux_52_i17_4_lut (.A(n7677[16]), .B(w_result[16]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i17_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i18_3_lut (.A(m_result[17]), .B(x_result[17]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i18_3_lut.init = 16'hcaca;
    LUT4 mux_52_i18_4_lut (.A(n7677[17]), .B(w_result[17]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i18_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i19_3_lut (.A(m_result[18]), .B(x_result[18]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i19_3_lut.init = 16'hcaca;
    LUT4 mux_52_i19_4_lut (.A(n7677[18]), .B(w_result[18]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i19_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i20_3_lut (.A(m_result[19]), .B(x_result[19]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i20_3_lut.init = 16'hcaca;
    LUT4 i14588_2_lut (.A(icache_refilling), .B(dcache_refilling), .Z(n19852)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14588_2_lut.init = 16'heeee;
    LUT4 i46_rep_22_4_lut (.A(n32128), .B(LM32D_CYC_O), .C(n32134), .D(n32132), 
         .Z(n30493)) /* synthesis lut_function=(A (B)+!A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1.v(400[8:19])
    defparam i46_rep_22_4_lut.init = 16'hc888;
    LUT4 mux_52_i20_4_lut (.A(n7677[19]), .B(w_result[19]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i20_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i21_3_lut (.A(m_result[20]), .B(x_result[20]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i21_3_lut.init = 16'hcaca;
    LUT4 mux_52_i21_4_lut (.A(n7677[20]), .B(w_result[20]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i21_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i22_3_lut (.A(m_result[21]), .B(x_result[21]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i22_3_lut.init = 16'hcaca;
    LUT4 mux_52_i22_4_lut (.A(n7677[21]), .B(w_result[21]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i22_4_lut.init = 16'hcac0;
    LUT4 i1_4_lut_adj_608 (.A(n33942), .B(n33944), .C(n33946), .D(n41283), 
         .Z(non_debug_exception_x)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1771[32] 1791[33])
    defparam i1_4_lut_adj_608.init = 16'heefe;
    LUT4 bypass_data_1_31__I_15_i23_3_lut (.A(m_result[22]), .B(x_result[22]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i23_3_lut.init = 16'hcaca;
    LUT4 mux_52_i23_4_lut (.A(n7677[22]), .B(w_result[22]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i23_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i24_3_lut (.A(m_result[23]), .B(x_result[23]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i24_3_lut.init = 16'hcaca;
    LUT4 mux_52_i24_4_lut (.A(n7677[23]), .B(w_result[23]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i24_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i25_3_lut (.A(m_result[24]), .B(x_result[24]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i25_3_lut.init = 16'hcaca;
    LUT4 mux_52_i25_4_lut (.A(n7677[24]), .B(w_result[24]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[24])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i25_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i26_3_lut (.A(m_result[25]), .B(x_result[25]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i26_3_lut.init = 16'hcaca;
    LUT4 mux_52_i26_4_lut (.A(n7677[25]), .B(w_result[25]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[25])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i26_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i27_3_lut (.A(m_result[26]), .B(x_result[26]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i27_3_lut.init = 16'hcaca;
    LUT4 mux_52_i27_4_lut (.A(n7677[26]), .B(w_result[26]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[26])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i27_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i28_3_lut (.A(m_result[27]), .B(x_result[27]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i28_3_lut.init = 16'hcaca;
    LUT4 mux_52_i28_4_lut (.A(n7677[27]), .B(w_result[27]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[27])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i28_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i29_3_lut (.A(m_result[28]), .B(x_result[28]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i29_3_lut.init = 16'hcaca;
    LUT4 mux_52_i29_4_lut (.A(n7677[28]), .B(w_result[28]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[28])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i29_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i30_3_lut (.A(m_result[29]), .B(x_result[29]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i30_3_lut.init = 16'hcaca;
    LUT4 mux_52_i30_4_lut (.A(n7677[29]), .B(w_result[29]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i30_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i31_3_lut (.A(m_result[30]), .B(x_result[30]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i31_3_lut.init = 16'hcaca;
    LUT4 mux_52_i31_4_lut (.A(n7677[30]), .B(w_result[30]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i31_4_lut.init = 16'hcac0;
    LUT4 bypass_data_1_31__I_15_i32_3_lut (.A(m_result[31]), .B(x_result[31]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_914[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_15_i32_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut (.A(store_m), .B(w_result_sel_load_x), .C(load_m), .Z(n32128)) /* synthesis lut_function=(A+(B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(365[5:16])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 mux_52_i32_4_lut (.A(n7677[31]), .B(w_result[31]), .C(raw_w_1), 
         .D(n6648), .Z(bypass_data_1_31__N_1044[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i32_4_lut.init = 16'hcac0;
    LUT4 mux_2953_i11_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7224), 
         .D(adder_result_x[12]), .Z(n7190[10])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2953_i11_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3055_i6_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra [5]), 
         .D(adder_result_x[7]), .Z(n7388[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3055_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3055_i3_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra [2]), 
         .D(adder_result_x[4]), .Z(n7388[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3055_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 n41751_bdd_3_lut (.A(n41751), .B(n41749), .C(x_result_sel_sext_x), 
         .Z(n41752)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41751_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_1099 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_431)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1099.init = 16'h0f0e;
    LUT4 n4_bdd_3_lut_34327 (.A(operand_w[14]), .B(multiplier_result_w[14]), 
         .C(w_result_sel_mul_w), .Z(n41142)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n4_bdd_3_lut_34327.init = 16'hcaca;
    LUT4 i14851_4_lut (.A(extended_immediate[31]), .B(n41179), .C(n41375), 
         .D(n41291), .Z(n2_adj_6196)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1558[5] 1563[12])
    defparam i14851_4_lut.init = 16'hc088;
    LUT4 i14852_4_lut (.A(extended_immediate[31]), .B(n41179), .C(n41374), 
         .D(n41291), .Z(n2_adj_6197)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1558[5] 1563[12])
    defparam i14852_4_lut.init = 16'hc088;
    LUT4 i14917_4_lut (.A(extended_immediate[31]), .B(n41179), .C(n41373), 
         .D(n41291), .Z(n2_adj_6198)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1558[5] 1563[12])
    defparam i14917_4_lut.init = 16'hc088;
    LUT4 i14926_4_lut (.A(extended_immediate[31]), .B(n41179), .C(n41372), 
         .D(n41291), .Z(n2_adj_6199)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1558[5] 1563[12])
    defparam i14926_4_lut.init = 16'hc088;
    LUT4 i14928_4_lut (.A(extended_immediate[31]), .B(n41179), .C(n41371), 
         .D(n41291), .Z(n2_adj_6200)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1558[5] 1563[12])
    defparam i14928_4_lut.init = 16'hc088;
    LUT4 i14931_4_lut (.A(extended_immediate[31]), .B(n41179), .C(n41370), 
         .D(n41291), .Z(n2_adj_6201)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1558[5] 1563[12])
    defparam i14931_4_lut.init = 16'hc088;
    LUT4 i14932_4_lut (.A(extended_immediate[31]), .B(n41179), .C(n41361), 
         .D(n41291), .Z(n2_adj_6202)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1558[5] 1563[12])
    defparam i14932_4_lut.init = 16'hc088;
    LUT4 i14933_4_lut (.A(extended_immediate[31]), .B(n41179), .C(n41369), 
         .D(n41291), .Z(n2_adj_6203)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1558[5] 1563[12])
    defparam i14933_4_lut.init = 16'hc088;
    LUT4 i14934_4_lut (.A(extended_immediate[31]), .B(n41179), .C(n41368), 
         .D(n41291), .Z(n2_adj_6204)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1558[5] 1563[12])
    defparam i14934_4_lut.init = 16'hc088;
    LUT4 mux_2953_i10_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7222), 
         .D(adder_result_x[11]), .Z(n7190[9])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2953_i10_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_rep_1100 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_430)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1100.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_1101 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_61)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1101.init = 16'h0f0e;
    LUT4 i1_4_lut_adj_609 (.A(n41291), .B(n41179), .C(n41348), .D(n41198), 
         .Z(n31335)) /* synthesis lut_function=(A (B (C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1558[5] 1563[12])
    defparam i1_4_lut_adj_609.init = 16'hc080;
    LUT4 i15252_4_lut (.A(extended_immediate[31]), .B(n41179), .C(n41377), 
         .D(n41291), .Z(n2_adj_6205)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1558[5] 1563[12])
    defparam i15252_4_lut.init = 16'hc088;
    LUT4 i1_2_lut_rep_1102 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_699)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1102.init = 16'h0f0e;
    LUT4 i15253_4_lut (.A(extended_immediate[31]), .B(n41179), .C(n41376), 
         .D(n41291), .Z(n2_adj_6206)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1558[5] 1563[12])
    defparam i15253_4_lut.init = 16'hc088;
    LUT4 i1_2_lut_rep_1103 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_700)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1103.init = 16'h0f0e;
    LUT4 mux_3055_i4_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra [3]), 
         .D(adder_result_x[5]), .Z(n7388[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3055_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_2953_i1_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7204), .D(adder_result_x[2]), 
         .Z(n7190[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2953_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_2953_i4_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7210), .D(adder_result_x[5]), 
         .Z(n7190[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2953_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_2953_i5_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7212), .D(adder_result_x[6]), 
         .Z(n7190[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2953_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_2953_i6_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7214), .D(adder_result_x[7]), 
         .Z(n7190[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2953_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_rep_1104 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_701)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1104.init = 16'h0f0e;
    LUT4 mux_2953_i7_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7216), .D(adder_result_x[8]), 
         .Z(n7190[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2953_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i12657_3_lut (.A(operand_m[0]), .B(condition_met_m), .C(m_result_sel_compare_m), 
         .Z(n17971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(443[5:25])
    defparam i12657_3_lut.init = 16'hcaca;
    LUT4 D_CYC_O_I_0_1_lut_rep_983 (.A(LM32D_CYC_O), .Z(n41388)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1789[8:27])
    defparam D_CYC_O_I_0_1_lut_rep_983.init = 16'h5555;
    LUT4 i2619_2_lut_2_lut_rep_984 (.A(LM32D_CYC_O), .B(dcache_refill_request), 
         .Z(n41389)) /* synthesis lut_function=(!(A+!(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1789[8:27])
    defparam i2619_2_lut_2_lut_rep_984.init = 16'h4444;
    LUT4 i7037_3_lut_4_lut_4_lut (.A(LM32D_CYC_O), .B(dcache_refill_request), 
         .C(n41217), .D(n41215), .Z(REF_CLK_c_enable_1234)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1789[8:27])
    defparam i7037_3_lut_4_lut_4_lut.init = 16'h5554;
    LUT4 mux_432_i1_3_lut (.A(branch_target_d[2]), .B(bypass_data_0[2]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i1_3_lut.init = 16'hcaca;
    LUT4 i12656_3_lut (.A(left_shift_result[31]), .B(left_shift_result[0]), 
         .C(direction_m), .Z(n17970)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(92[5:16])
    defparam i12656_3_lut.init = 16'hcaca;
    LUT4 mux_3055_i11_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra [10]), 
         .D(adder_result_x[12]), .Z(n7388[10])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3055_i11_3_lut_4_lut.init = 16'hf4b0;
    CCU2C operand_0_x_31__I_0_27 (.A0(operand_1_x[13]), .B0(operand_0_x[13]), 
          .C0(operand_1_x[12]), .D0(operand_0_x[12]), .A1(operand_1_x[11]), 
          .B1(operand_0_x[11]), .C1(operand_1_x[10]), .D1(operand_0_x[10]), 
          .CIN(n27362), .COUT(n27363));
    defparam operand_0_x_31__I_0_27.INIT0 = 16'h9009;
    defparam operand_0_x_31__I_0_27.INIT1 = 16'h9009;
    defparam operand_0_x_31__I_0_27.INJECT1_0 = "YES";
    defparam operand_0_x_31__I_0_27.INJECT1_1 = "YES";
    LUT4 mux_3055_i10_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra [9]), 
         .D(adder_result_x[11]), .Z(n7388[9])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3055_i10_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3055_i9_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra [8]), 
         .D(adder_result_x[10]), .Z(n7388[8])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3055_i9_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3055_i8_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra [7]), 
         .D(adder_result_x[9]), .Z(n7388[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3055_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_2953_i8_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7218), .D(adder_result_x[9]), 
         .Z(n7190[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2953_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3115_i9_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra_adj_6257 [8]), 
         .D(adder_result_x[12]), .Z(n7502[8])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3115_i9_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3115_i8_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra_adj_6257 [7]), 
         .D(adder_result_x[11]), .Z(n7502[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3115_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3115_i7_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra_adj_6257 [6]), 
         .D(adder_result_x[10]), .Z(n7502[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3115_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3115_i6_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra_adj_6257 [5]), 
         .D(adder_result_x[9]), .Z(n7502[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3115_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3115_i5_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra_adj_6257 [4]), 
         .D(adder_result_x[8]), .Z(n7502[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3115_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_4_lut_adj_610 (.A(n41232), .B(REF_CLK_c_enable_388), .C(n41233), 
         .D(n34898), .Z(eba_31__N_1111)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_610.init = 16'h0800;
    LUT4 mux_3115_i4_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra_adj_6257 [3]), 
         .D(adder_result_x[7]), .Z(n7502[3])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3115_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3115_i3_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra_adj_6257 [2]), 
         .D(adder_result_x[6]), .Z(n7502[2])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3115_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3115_i2_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra_adj_6257 [1]), 
         .D(adder_result_x[5]), .Z(n7502[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3115_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3115_i1_3_lut_4_lut (.A(n41233), .B(n41232), .C(\genblk1.ra_adj_6257 [0]), 
         .D(adder_result_x[4]), .Z(n7502[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_3115_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_2987_i11_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7290), 
         .D(adder_result_x[12]), .Z(n7256[10])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2987_i11_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_2987_i10_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7288), 
         .D(adder_result_x[11]), .Z(n7256[9])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2987_i10_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_2987_i9_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7286), .D(adder_result_x[10]), 
         .Z(n7256[8])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2987_i9_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_2987_i8_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7284), .D(adder_result_x[9]), 
         .Z(n7256[7])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2987_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_2987_i7_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7282), .D(adder_result_x[8]), 
         .Z(n7256[6])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2987_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_2987_i6_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7280), .D(adder_result_x[7]), 
         .Z(n7256[5])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2987_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_2987_i5_3_lut_4_lut (.A(n41233), .B(n41232), .C(n7278), .D(adder_result_x[6]), 
         .Z(n7256[4])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam mux_2987_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_adj_611 (.A(exception_m), .B(n17972), .Z(operand_w_31__N_850[0])) /* synthesis lut_function=(!(A+!(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i1_2_lut_adj_611.init = 16'h4444;
    LUT4 i1_2_lut_rep_1073 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_716)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1073.init = 16'h0f0e;
    LUT4 i1_2_lut_3_lut_4_lut (.A(cycles_5__N_2934), .B(n41231), .C(n41350), 
         .D(n41233), .Z(n32264)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i1_2_lut_rep_1074 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_717)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1074.init = 16'h0f0e;
    LUT4 i1_4_lut_adj_612 (.A(n41360), .B(n45171), .C(data_bus_error_exception), 
         .D(n9308), .Z(memop_pc_w_31__N_1229)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2618[16] 2622[17])
    defparam i1_4_lut_adj_612.init = 16'h0800;
    LUT4 load_q_m_I_0_2_lut (.A(load_m), .B(store_m), .Z(n9308)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2620[16] 2622[17])
    defparam load_q_m_I_0_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_rep_778_3_lut_4_lut (.A(cycles_5__N_2934), .B(n41231), 
         .C(REF_CLK_c_enable_388), .D(n41233), .Z(n41183)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i1_2_lut_rep_778_3_lut_4_lut.init = 16'h00e0;
    LUT4 i1_3_lut_4_lut_3_lut (.A(cycles_5__N_2934), .B(n41201), .C(n41233), 
         .Z(n32608)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i1_3_lut_4_lut_3_lut.init = 16'h0202;
    LUT4 i1_3_lut_4_lut_adj_613 (.A(cycles_5__N_2934), .B(n41231), .C(n41233), 
         .D(x_result_sel_csr_d), .Z(n19987)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;
    defparam i1_3_lut_4_lut_adj_613.init = 16'hf1ff;
    LUT4 i14594_3_lut (.A(write_idx_x[0]), .B(non_debug_exception_x), .C(n41417), 
         .Z(write_idx_m_4__N_1162[0])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2532[18] 2535[47])
    defparam i14594_3_lut.init = 16'h3232;
    LUT4 i15308_2_lut_3_lut (.A(n41417), .B(non_debug_exception_x), .C(write_idx_x[1]), 
         .Z(write_idx_m_4__N_1162[1])) /* synthesis lut_function=(A+(B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2532[18] 2535[47])
    defparam i15308_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_1075 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_718)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1075.init = 16'h0f0e;
    LUT4 n4_bdd_3_lut_34332 (.A(operand_w[13]), .B(multiplier_result_w[13]), 
         .C(w_result_sel_mul_w), .Z(n41146)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n4_bdd_3_lut_34332.init = 16'hcaca;
    LUT4 i15310_2_lut_3_lut (.A(n41417), .B(non_debug_exception_x), .C(write_idx_x[3]), 
         .Z(write_idx_m_4__N_1162[3])) /* synthesis lut_function=(A+(B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2532[18] 2535[47])
    defparam i15310_2_lut_3_lut.init = 16'hfefe;
    LUT4 i15311_2_lut_3_lut (.A(n41417), .B(non_debug_exception_x), .C(write_idx_x[4]), 
         .Z(write_idx_m_4__N_1162[4])) /* synthesis lut_function=(A+(B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2532[18] 2535[47])
    defparam i15311_2_lut_3_lut.init = 16'hfefe;
    LUT4 i15309_2_lut_3_lut (.A(n41417), .B(non_debug_exception_x), .C(write_idx_x[2]), 
         .Z(write_idx_m_4__N_1162[2])) /* synthesis lut_function=(A+(B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2532[18] 2535[47])
    defparam i15309_2_lut_3_lut.init = 16'hfefe;
    FD1P3DX valid_d_663 (.D(n31132), .SP(REF_CLK_c_enable_1622), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(valid_d)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2264[5] 2299[8])
    defparam valid_d_663.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_1076 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_719)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1076.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_1077 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_720)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1077.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_1078 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_721)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1078.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_1079 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_722)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1079.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_1080 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_723)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1080.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_1081 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_724)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1081.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_1082 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_725)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1082.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_1083 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_726)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1083.init = 16'h0f0e;
    LUT4 i1_4_lut_adj_614 (.A(n35639), .B(dcache_refill_request), .C(n35022), 
         .D(operand_1_x[0]), .Z(n34986)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_614.init = 16'h1000;
    LUT4 i1_3_lut_adj_615 (.A(dcache_refill_request), .B(valid_x), .C(bret_x), 
         .Z(n35030)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut_adj_615.init = 16'h4040;
    LUT4 i1_2_lut_adj_616 (.A(valid_x), .B(csr_write_enable_x), .Z(n35022)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_616.init = 16'h8888;
    LUT4 i1_4_lut_adj_617 (.A(n41232), .B(n41202), .C(n45068), .D(n41233), 
         .Z(n31804)) /* synthesis lut_function=(A (B (C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i1_4_lut_adj_617.init = 16'hc080;
    LUT4 i1_2_lut_rep_1084 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_727)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1084.init = 16'h0f0e;
    LUT4 n10760_bdd_3_lut_33750_3_lut (.A(csr_x[0]), .B(eba[11]), .C(csr_x[3]), 
         .Z(n39323)) /* synthesis lut_function=(!(A ((C)+!B)+!A (C))) */ ;
    defparam n10760_bdd_3_lut_33750_3_lut.init = 16'h0d0d;
    LUT4 mux_2223_i1_4_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(jrx_csr_read_data[0]), 
         .Z(n5780[0])) /* synthesis lut_function=(A (B (C))+!A !(B)) */ ;
    defparam mux_2223_i1_4_lut_3_lut.init = 16'h9191;
    LUT4 mux_2223_i2_4_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(jrx_csr_read_data[1]), 
         .Z(n5780[1])) /* synthesis lut_function=(A (B (C))+!A !(B)) */ ;
    defparam mux_2223_i2_4_lut_3_lut.init = 16'h9191;
    LUT4 mux_2223_i3_4_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(jrx_csr_read_data[2]), 
         .Z(n5780[2])) /* synthesis lut_function=(A (B (C))+!A !(B)) */ ;
    defparam mux_2223_i3_4_lut_3_lut.init = 16'h9191;
    LUT4 i14062_3_lut (.A(operand_m[25]), .B(dcache_refill_address[25]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(676[6:27])
    defparam i14062_3_lut.init = 16'hcaca;
    LUT4 eba_8__bdd_4_lut_4_lut (.A(csr_x[0]), .B(csr_x[3]), .C(n39310), 
         .D(eba[8]), .Z(n41168)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;
    defparam eba_8__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 mux_2223_i4_4_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(jrx_csr_read_data[3]), 
         .Z(n5780[3])) /* synthesis lut_function=(A (B (C))+!A !(B)) */ ;
    defparam mux_2223_i4_4_lut_3_lut.init = 16'h9191;
    LUT4 mux_2223_i7_4_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(jrx_csr_read_data[6]), 
         .Z(n5780[6])) /* synthesis lut_function=(A (B (C))+!A !(B)) */ ;
    defparam mux_2223_i7_4_lut_3_lut.init = 16'h9191;
    LUT4 i14047_3_lut (.A(operand_m[27]), .B(dcache_refill_address[27]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(676[6:27])
    defparam i14047_3_lut.init = 16'hcaca;
    LUT4 mux_2223_i8_4_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(jrx_csr_read_data[7]), 
         .Z(n5780[7])) /* synthesis lut_function=(A (B (C))+!A !(B)) */ ;
    defparam mux_2223_i8_4_lut_3_lut.init = 16'h9191;
    LUT4 i1_2_lut_rep_1105 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_702)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1105.init = 16'h0f0e;
    LUT4 n4_bdd_3_lut_34337 (.A(operand_w[12]), .B(multiplier_result_w[12]), 
         .C(w_result_sel_mul_w), .Z(n41150)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n4_bdd_3_lut_34337.init = 16'hcaca;
    LUT4 i1_4_lut_adj_618 (.A(n41196), .B(n45175), .C(branch_taken_m), 
         .D(n32630), .Z(n32636)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_618.init = 16'h0400;
    LUT4 i1_4_lut_adj_619 (.A(n41216), .B(n41435), .C(cycles_5__N_2934), 
         .D(valid_d), .Z(n32630)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_619.init = 16'h1000;
    LUT4 n4_bdd_3_lut_34342 (.A(operand_w[11]), .B(multiplier_result_w[11]), 
         .C(w_result_sel_mul_w), .Z(n41154)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n4_bdd_3_lut_34342.init = 16'hcaca;
    LUT4 i1_2_lut_rep_1106 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_703)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1106.init = 16'h0f0e;
    LUT4 i4039_2_lut_rep_986 (.A(csr_x[3]), .B(csr_x[0]), .Z(n41391)) /* synthesis lut_function=(A (B)) */ ;
    defparam i4039_2_lut_rep_986.init = 16'h8888;
    LUT4 n4_bdd_3_lut_34347 (.A(operand_w[10]), .B(multiplier_result_w[10]), 
         .C(w_result_sel_mul_w), .Z(n41158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n4_bdd_3_lut_34347.init = 16'hcaca;
    LUT4 i1_3_lut_rep_768_4_lut (.A(n41232), .B(n41233), .C(n15), .D(n41196), 
         .Z(REF_CLK_c_enable_1425)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_3_lut_rep_768_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(csr_x[3]), .B(csr_x[0]), .C(im[7]), 
         .D(n41308), .Z(n19)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_3_lut_4_lut_adj_620 (.A(n41417), .B(non_debug_exception_x), 
         .C(w_result_sel_mul_x), .D(n45171), .Z(n12394)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam i1_2_lut_3_lut_4_lut_adj_620.init = 16'h10f0;
    LUT4 i14597_2_lut_3_lut (.A(n41417), .B(non_debug_exception_x), .C(write_enable_x), 
         .Z(write_enable_m_N_1339)) /* synthesis lut_function=(A+(B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam i14597_2_lut_3_lut.init = 16'hfefe;
    LUT4 i14596_2_lut_3_lut (.A(n41417), .B(non_debug_exception_x), .C(branch_target_x[2]), 
         .Z(branch_target_m_31__N_1167[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam i14596_2_lut_3_lut.init = 16'h1010;
    FD1S3DX write_idx_w_i0_rep_1069 (.D(write_idx_m[0]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n45103)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_w_i0_rep_1069.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut_adj_621 (.A(n7_adj_6195), .B(n41420), .C(n30493), 
         .D(n41436), .Z(n30089)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_621.init = 16'h0400;
    LUT4 mux_1680_i24_3_lut_4_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[15]), 
         .D(operand_0_x[7]), .Z(sext_result_x[31])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1576[24:49])
    defparam mux_1680_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_622 (.A(csr_x[3]), .B(csr_x[0]), 
         .C(im[3]), .D(n41308), .Z(n17)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_622.init = 16'h0040;
    LUT4 i1_2_lut_3_lut_4_lut_adj_623 (.A(n41417), .B(non_debug_exception_x), 
         .C(w_result_sel_load_x), .D(n45171), .Z(n12410)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam i1_2_lut_3_lut_4_lut_adj_623.init = 16'h10f0;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_624 (.A(csr_x[3]), .B(csr_x[0]), 
         .C(im[6]), .D(n41308), .Z(n18)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_624.init = 16'h0040;
    LUT4 n4_bdd_3_lut_34352 (.A(operand_w[9]), .B(multiplier_result_w[9]), 
         .C(w_result_sel_mul_w), .Z(n41162)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n4_bdd_3_lut_34352.init = 16'hcaca;
    LUT4 i1_2_lut_rep_1107 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_704)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1107.init = 16'h0f0e;
    FD1P3DX x_result_sel_add_x_675 (.D(n31549), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(x_result_sel_add_x)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam x_result_sel_add_x_675.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_1108 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_705)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1108.init = 16'h0f0e;
    LUT4 i15066_2_lut_3_lut (.A(n41417), .B(non_debug_exception_x), .C(branch_target_x[3]), 
         .Z(branch_target_m_31__N_1167[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam i15066_2_lut_3_lut.init = 16'h1010;
    LUT4 i15067_2_lut_3_lut (.A(n41417), .B(non_debug_exception_x), .C(branch_target_x[4]), 
         .Z(branch_target_m_31__N_1167[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam i15067_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_4_lut_adj_625 (.A(n20581), .B(REF_CLK_c_enable_388), .C(n41232), 
         .D(n34880), .Z(REF_CLK_c_enable_1335)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_625.init = 16'h4000;
    LUT4 i1_4_lut_adj_626 (.A(n41233), .B(n41313), .C(n34874), .D(REF_CLK_c_enable_391), 
         .Z(n34880)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_626.init = 16'h1000;
    LUT4 mux_508_i5_4_lut_4_lut (.A(n41417), .B(non_debug_exception_x), 
         .C(n35412), .D(branch_target_x[6]), .Z(branch_target_m_31__N_1167[4])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i5_4_lut_4_lut.init = 16'h5140;
    FD1S3DX write_idx_w_i1_rep_1065 (.D(write_idx_m[1]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n45099)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_w_i1_rep_1065.GSR = "ENABLED";
    LUT4 i33078_2_lut_rep_994 (.A(non_debug_exception_w), .B(valid_w), .Z(REF_CLK_c_enable_391)) /* synthesis lut_function=(!(A (B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2008[34:90])
    defparam i33078_2_lut_rep_994.init = 16'h7777;
    LUT4 n41753_bdd_3_lut (.A(n41753), .B(adder_result_x[11]), .C(x_result_sel_add_x), 
         .Z(x_result[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41753_bdd_3_lut.init = 16'hcaca;
    LUT4 logic_result_x_12__bdd_4_lut_34522 (.A(n39327), .B(n5915), .C(n39326), 
         .D(csr_x[2]), .Z(n41755)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam logic_result_x_12__bdd_4_lut_34522.init = 16'hc088;
    LUT4 i1_2_lut_rep_1109 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_706)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1109.init = 16'h0f0e;
    LUT4 i4107_3_lut_4_lut (.A(non_debug_exception_w), .B(valid_w), .C(ie), 
         .D(\operand_1_x[1] ), .Z(n9401)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2008[34:90])
    defparam i4107_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_627 (.A(n41317), .B(REF_CLK_c_enable_388), .C(n41394), 
         .D(n41233), .Z(n31501)) /* synthesis lut_function=(!((B (C)+!B (C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_627.init = 16'h0a08;
    LUT4 i4012_3_lut (.A(valid_w), .B(debug_exception_w), .C(non_debug_exception_w), 
         .Z(jtag_reg_d_7__N_515)) /* synthesis lut_function=(A (B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1184[30:76])
    defparam i4012_3_lut.init = 16'ha8a8;
    LUT4 logic_result_x_12__bdd_4_lut_35512 (.A(size_x[1]), .B(size_x[0]), 
         .C(operand_0_x[12]), .D(operand_0_x[7]), .Z(n41756)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam logic_result_x_12__bdd_4_lut_35512.init = 16'hf1e0;
    LUT4 logic_result_x_12__bdd_3_lut_35513 (.A(size_x[1]), .B(size_x[0]), 
         .C(operand_0_x[12]), .Z(n41757)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam logic_result_x_12__bdd_3_lut_35513.init = 16'hacac;
    LUT4 n4_bdd_3_lut (.A(operand_w[8]), .B(multiplier_result_w[8]), .C(w_result_sel_mul_w), 
         .Z(n41166)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n4_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_628 (.A(n41232), .B(n41233), .C(n41448), .D(n41393), 
         .Z(n33932)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam i1_4_lut_adj_628.init = 16'hfffd;
    LUT4 i1_2_lut_rep_1085 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_728)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1085.init = 16'h0f0e;
    LUT4 debug_exception_w_I_0_2_lut_rep_996 (.A(debug_exception_w), .B(valid_w), 
         .Z(n41401)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2007[30:82])
    defparam debug_exception_w_I_0_2_lut_rep_996.init = 16'h8888;
    LUT4 n41758_bdd_3_lut (.A(n41758), .B(n41756), .C(x_result_sel_sext_x), 
         .Z(n41759)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41758_bdd_3_lut.init = 16'hcaca;
    LUT4 bie_I_134_3_lut_4_lut (.A(debug_exception_w), .B(valid_w), .C(ie), 
         .D(operand_1_x[2]), .Z(bie_N_3274)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2007[30:82])
    defparam bie_I_134_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_1110 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_707)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1110.init = 16'h0f0e;
    LUT4 i1_4_lut_adj_629 (.A(branch_flushX_m), .B(n41233), .C(n41240), 
         .D(n34936), .Z(n34942)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam i1_4_lut_adj_629.init = 16'hfffe;
    LUT4 i1_4_lut_adj_630 (.A(n35767), .B(n11934), .C(csr_write_enable_x), 
         .D(dcache_refill_request), .Z(n34936)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1907[21] 1911[22])
    defparam i1_4_lut_adj_630.init = 16'hffdf;
    LUT4 i30606_2_lut (.A(\operand_1_x[1] ), .B(valid_x), .Z(n35767)) /* synthesis lut_function=(A (B)) */ ;
    defparam i30606_2_lut.init = 16'h8888;
    CCU2C operand_0_x_31__I_0_25 (.A0(operand_1_x[17]), .B0(operand_0_x[17]), 
          .C0(operand_1_x[16]), .D0(operand_0_x[16]), .A1(operand_1_x[15]), 
          .B1(operand_0_x[15]), .C1(operand_1_x[14]), .D1(operand_0_x[14]), 
          .CIN(n27361), .COUT(n27362));
    defparam operand_0_x_31__I_0_25.INIT0 = 16'h9009;
    defparam operand_0_x_31__I_0_25.INIT1 = 16'h9009;
    defparam operand_0_x_31__I_0_25.INJECT1_0 = "YES";
    defparam operand_0_x_31__I_0_25.INJECT1_1 = "YES";
    LUT4 size_x_1__I_0_743_i3_2_lut_rep_997 (.A(size_x[0]), .B(size_x[1]), 
         .Z(n41402)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1576[24:49])
    defparam size_x_1__I_0_743_i3_2_lut_rep_997.init = 16'heeee;
    CCU2C operand_0_x_31__I_0_23 (.A0(operand_1_x[21]), .B0(operand_0_x[21]), 
          .C0(operand_1_x[20]), .D0(operand_0_x[20]), .A1(operand_1_x[19]), 
          .B1(operand_0_x[19]), .C1(operand_1_x[18]), .D1(operand_0_x[18]), 
          .CIN(n27360), .COUT(n27361));
    defparam operand_0_x_31__I_0_23.INIT0 = 16'h9009;
    defparam operand_0_x_31__I_0_23.INIT1 = 16'h9009;
    defparam operand_0_x_31__I_0_23.INJECT1_0 = "YES";
    defparam operand_0_x_31__I_0_23.INJECT1_1 = "YES";
    LUT4 i1_3_lut_rep_1048 (.A(dcache_refill_request), .B(branch_flushX_m), 
         .C(valid_x), .Z(n45068)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_3_lut_rep_1048.init = 16'h1010;
    CCU2C operand_0_x_31__I_0_21 (.A0(operand_1_x[25]), .B0(operand_0_x[25]), 
          .C0(operand_1_x[24]), .D0(operand_0_x[24]), .A1(operand_1_x[23]), 
          .B1(operand_0_x[23]), .C1(operand_1_x[22]), .D1(operand_0_x[22]), 
          .CIN(n27359), .COUT(n27360));
    defparam operand_0_x_31__I_0_21.INIT0 = 16'h9009;
    defparam operand_0_x_31__I_0_21.INIT1 = 16'h9009;
    defparam operand_0_x_31__I_0_21.INJECT1_0 = "YES";
    defparam operand_0_x_31__I_0_21.INJECT1_1 = "YES";
    LUT4 i1_2_lut_rep_1087 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_443)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1087.init = 16'h0f0e;
    LUT4 n41760_bdd_3_lut (.A(n41760), .B(adder_result_x[12]), .C(x_result_sel_add_x), 
         .Z(x_result[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41760_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_1111 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_708)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1111.init = 16'h0f0e;
    LUT4 logic_result_x_13__bdd_4_lut_34527 (.A(n39330), .B(n5915), .C(n39329), 
         .D(csr_x[2]), .Z(n41762)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam logic_result_x_13__bdd_4_lut_34527.init = 16'hc088;
    LUT4 i1_2_lut_rep_1112 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_709)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1112.init = 16'h0f0e;
    LUT4 logic_result_x_13__bdd_4_lut_35331 (.A(size_x[1]), .B(size_x[0]), 
         .C(operand_0_x[13]), .D(operand_0_x[7]), .Z(n41763)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam logic_result_x_13__bdd_4_lut_35331.init = 16'hf1e0;
    LUT4 logic_result_x_13__bdd_3_lut_35332 (.A(size_x[1]), .B(size_x[0]), 
         .C(operand_0_x[13]), .Z(n41764)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam logic_result_x_13__bdd_3_lut_35332.init = 16'hacac;
    LUT4 i1_2_lut_rep_1113 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_710)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1113.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_1114 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_711)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1114.init = 16'h0f0e;
    LUT4 bypass_data_0_31__I_0_i32_3_lut (.A(bypass_data_0[31]), .B(pc_f[31]), 
         .C(n41208), .Z(d_result_0[31])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i32_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i31_3_lut (.A(bypass_data_0[30]), .B(pc_f[30]), 
         .C(n41208), .Z(d_result_0[30])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i31_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i30_3_lut (.A(bypass_data_0[29]), .B(pc_f[29]), 
         .C(n41208), .Z(d_result_0[29])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i30_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i29_3_lut (.A(bypass_data_0[28]), .B(pc_f[28]), 
         .C(n41208), .Z(d_result_0[28])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i29_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i28_3_lut (.A(bypass_data_0[27]), .B(pc_f[27]), 
         .C(n41208), .Z(d_result_0[27])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i28_3_lut.init = 16'hacac;
    CCU2C operand_0_x_31__I_0_19 (.A0(operand_1_x[29]), .B0(operand_0_x[29]), 
          .C0(operand_1_x[28]), .D0(operand_0_x[28]), .A1(operand_1_x[27]), 
          .B1(operand_0_x[27]), .C1(operand_1_x[26]), .D1(operand_0_x[26]), 
          .CIN(n27358), .COUT(n27359));
    defparam operand_0_x_31__I_0_19.INIT0 = 16'h9009;
    defparam operand_0_x_31__I_0_19.INIT1 = 16'h9009;
    defparam operand_0_x_31__I_0_19.INJECT1_0 = "YES";
    defparam operand_0_x_31__I_0_19.INJECT1_1 = "YES";
    LUT4 bypass_data_0_31__I_0_i27_3_lut (.A(bypass_data_0[26]), .B(pc_f[26]), 
         .C(n41208), .Z(d_result_0[26])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i27_3_lut.init = 16'hacac;
    CCU2C operand_0_x_31__I_0_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(operand_1_x[31]), .B1(operand_0_x[31]), .C1(operand_1_x[30]), 
          .D1(operand_0_x[30]), .COUT(n27358));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1585[19:45])
    defparam operand_0_x_31__I_0_0.INIT0 = 16'h000F;
    defparam operand_0_x_31__I_0_0.INIT1 = 16'h9009;
    defparam operand_0_x_31__I_0_0.INJECT1_0 = "NO";
    defparam operand_0_x_31__I_0_0.INJECT1_1 = "YES";
    LUT4 bypass_data_0_31__I_0_i26_3_lut (.A(bypass_data_0[25]), .B(pc_f[25]), 
         .C(n41208), .Z(d_result_0[25])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i26_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i25_3_lut (.A(bypass_data_0[24]), .B(pc_f[24]), 
         .C(n41208), .Z(d_result_0[24])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i25_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i24_3_lut (.A(bypass_data_0[23]), .B(pc_f[23]), 
         .C(n41208), .Z(d_result_0[23])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i24_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i23_3_lut (.A(bypass_data_0[22]), .B(pc_f[22]), 
         .C(n41208), .Z(d_result_0[22])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i23_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i22_3_lut (.A(bypass_data_0[21]), .B(pc_f[21]), 
         .C(n41208), .Z(d_result_0[21])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i22_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i21_3_lut (.A(bypass_data_0[20]), .B(pc_f[20]), 
         .C(n41208), .Z(d_result_0[20])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i21_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i20_3_lut (.A(bypass_data_0[19]), .B(pc_f[19]), 
         .C(n41208), .Z(d_result_0[19])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i20_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i19_3_lut (.A(bypass_data_0[18]), .B(pc_f[18]), 
         .C(n41208), .Z(d_result_0[18])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i19_3_lut.init = 16'hacac;
    LUT4 n41765_bdd_3_lut (.A(n41765), .B(n41763), .C(x_result_sel_sext_x), 
         .Z(n41766)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41765_bdd_3_lut.init = 16'hcaca;
    LUT4 bypass_data_0_31__I_0_i18_3_lut (.A(bypass_data_0[17]), .B(pc_f[17]), 
         .C(n41208), .Z(d_result_0[17])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i18_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i17_3_lut (.A(bypass_data_0[16]), .B(pc_f[16]), 
         .C(n41208), .Z(d_result_0[16])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i17_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i16_3_lut (.A(bypass_data_0[15]), .B(pc_f[15]), 
         .C(n41208), .Z(d_result_0[15])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i16_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i15_3_lut (.A(bypass_data_0[14]), .B(pc_f[14]), 
         .C(n41208), .Z(d_result_0[14])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i15_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i14_3_lut (.A(bypass_data_0[13]), .B(pc_f[13]), 
         .C(n41208), .Z(d_result_0[13])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i14_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i13_3_lut (.A(bypass_data_0[12]), .B(pc_f[12]), 
         .C(n41208), .Z(d_result_0[12])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i13_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i12_3_lut (.A(bypass_data_0[11]), .B(pc_f[11]), 
         .C(n41208), .Z(d_result_0[11])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i12_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_rep_1008 (.A(csr_x[0]), .B(csr_x[1]), .Z(n41413)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_1008.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_631 (.A(csr_x[0]), .B(csr_x[1]), .C(n41448), 
         .D(n41233), .Z(n34464)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_3_lut_4_lut_adj_631.init = 16'hfff7;
    LUT4 i1_2_lut_rep_1009 (.A(data_bus_error_exception), .B(reset_exception), 
         .Z(n41414)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1771[32] 1791[33])
    defparam i1_2_lut_rep_1009.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_632 (.A(data_bus_error_exception), .B(reset_exception), 
         .C(valid_x), .D(scall_x), .Z(n33944)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1771[32] 1791[33])
    defparam i1_3_lut_4_lut_adj_632.init = 16'hfeee;
    LUT4 i1_3_lut_4_lut_adj_633 (.A(data_bus_error_exception), .B(reset_exception), 
         .C(n41415), .D(divide_by_zero_x), .Z(n35412)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1771[32] 1791[33])
    defparam i1_3_lut_4_lut_adj_633.init = 16'h1011;
    LUT4 bus_error_x_I_0_2_lut_rep_1010 (.A(bus_error_x), .B(valid_x), .Z(n41415)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1750[42] 1752[43])
    defparam bus_error_x_I_0_2_lut_rep_1010.init = 16'h8888;
    LUT4 i15034_3_lut_4_lut (.A(bus_error_x), .B(valid_x), .C(n41417), 
         .D(data_bus_error_exception), .Z(eid_x_2__N_1009[2])) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A ((D)+!C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1750[42] 1752[43])
    defparam i15034_3_lut_4_lut.init = 16'hff07;
    LUT4 i1_2_lut_3_lut_adj_634 (.A(bus_error_x), .B(valid_x), .C(divide_by_zero_x), 
         .Z(n33942)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1750[42] 1752[43])
    defparam i1_2_lut_3_lut_adj_634.init = 16'hf8f8;
    LUT4 bypass_data_0_31__I_0_i11_3_lut (.A(bypass_data_0[10]), .B(pc_f[10]), 
         .C(n41208), .Z(d_result_0[10])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i11_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i10_3_lut (.A(bypass_data_0[9]), .B(pc_f[9]), 
         .C(n41208), .Z(d_result_0[9])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i10_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i9_3_lut (.A(bypass_data_0[8]), .B(pc_f[8]), 
         .C(n41208), .Z(d_result_0[8])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i9_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i8_3_lut (.A(bypass_data_0[7]), .B(pc_f[7]), 
         .C(n41208), .Z(d_result_0[7])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i8_3_lut.init = 16'hacac;
    PFUMX i34535 (.BLUT(n41776), .ALUT(n41772), .C0(x_result_sel_csr_x), 
          .Z(n41777));
    LUT4 bypass_data_0_31__I_0_i7_3_lut (.A(bypass_data_0[6]), .B(pc_f[6]), 
         .C(n41208), .Z(d_result_0[6])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i7_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i6_3_lut (.A(bypass_data_0[5]), .B(pc_f[5]), 
         .C(n41208), .Z(d_result_0[5])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i6_3_lut.init = 16'hacac;
    LUT4 breakpoint_exception_I_65_3_lut_rep_1012 (.A(break_x), .B(jtag_break), 
         .C(valid_x), .Z(n41417)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam breakpoint_exception_I_65_3_lut_rep_1012.init = 16'hecec;
    LUT4 bypass_data_0_31__I_0_i5_3_lut (.A(bypass_data_0[4]), .B(pc_f[4]), 
         .C(n41208), .Z(d_result_0[4])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i5_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i4_3_lut (.A(bypass_data_0[3]), .B(pc_f[3]), 
         .C(n41208), .Z(d_result_0[3])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i4_3_lut.init = 16'hacac;
    LUT4 bypass_data_0_31__I_0_i3_3_lut (.A(bypass_data_0[2]), .B(pc_f[2]), 
         .C(n41208), .Z(d_result_0[2])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1557[18:69])
    defparam bypass_data_0_31__I_0_i3_3_lut.init = 16'hacac;
    LUT4 debug_exception_x_I_0_2_lut_rep_797_4_lut (.A(break_x), .B(jtag_break), 
         .C(valid_x), .D(non_debug_exception_x), .Z(n41202)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam debug_exception_x_I_0_2_lut_rep_797_4_lut.init = 16'hffec;
    LUT4 n41767_bdd_3_lut (.A(n41767), .B(adder_result_x[13]), .C(x_result_sel_add_x), 
         .Z(x_result[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41767_bdd_3_lut.init = 16'hcaca;
    LUT4 logic_result_x_14__bdd_3_lut_35124 (.A(size_x[1]), .B(size_x[0]), 
         .C(operand_0_x[14]), .Z(n41774)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam logic_result_x_14__bdd_3_lut_35124.init = 16'hacac;
    LUT4 logic_result_x_14__bdd_4_lut_35123 (.A(size_x[1]), .B(size_x[0]), 
         .C(operand_0_x[14]), .D(operand_0_x[7]), .Z(n41773)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam logic_result_x_14__bdd_4_lut_35123.init = 16'hf1e0;
    LUT4 logic_result_x_14__bdd_4_lut_34532 (.A(n39333), .B(n5915), .C(n39332), 
         .D(csr_x[2]), .Z(n41772)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam logic_result_x_14__bdd_4_lut_34532.init = 16'hc088;
    LUT4 i1_2_lut_rep_1015 (.A(state[2]), .B(state_adj_6256[1]), .Z(n41420)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_1015.init = 16'h8888;
    LUT4 i1_3_lut_rep_828_4_lut (.A(state[2]), .B(state_adj_6256[1]), .C(n7_adj_6195), 
         .D(n30493), .Z(n41233)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_3_lut_rep_828_4_lut.init = 16'hfff7;
    LUT4 mux_432_i2_3_lut (.A(branch_target_d[3]), .B(bypass_data_0[3]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i2_3_lut.init = 16'hcaca;
    LUT4 mux_432_i3_3_lut (.A(branch_target_d[4]), .B(bypass_data_0[4]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i3_3_lut.init = 16'hcaca;
    LUT4 mux_432_i4_3_lut (.A(branch_target_d[5]), .B(bypass_data_0[5]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i4_3_lut.init = 16'hcaca;
    LUT4 mux_432_i5_3_lut (.A(branch_target_d[6]), .B(bypass_data_0[6]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i5_3_lut.init = 16'hcaca;
    LUT4 mux_432_i6_3_lut (.A(branch_target_d[7]), .B(bypass_data_0[7]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i6_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_rep_844_4_lut (.A(state[2]), .B(state_adj_6256[1]), .C(n30493), 
         .D(n7_adj_6195), .Z(REF_CLK_c_enable_1304)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_rep_844_4_lut.init = 16'h0008;
    PFUMX i34533 (.BLUT(logic_result_x[14]), .ALUT(n41774), .C0(n36757), 
          .Z(n41775));
    LUT4 mux_432_i7_3_lut (.A(branch_target_d[8]), .B(bypass_data_0[8]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i7_3_lut.init = 16'hcaca;
    LUT4 mux_432_i8_3_lut (.A(branch_target_d[9]), .B(bypass_data_0[9]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i8_3_lut.init = 16'hcaca;
    LUT4 mux_432_i9_3_lut (.A(branch_target_d[10]), .B(bypass_data_0[10]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i9_3_lut.init = 16'hcaca;
    LUT4 mux_432_i10_3_lut (.A(branch_target_d[11]), .B(bypass_data_0[11]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i10_3_lut.init = 16'hcaca;
    LUT4 mux_432_i11_3_lut (.A(branch_target_d[12]), .B(bypass_data_0[12]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i11_3_lut.init = 16'hcaca;
    LUT4 mux_432_i12_3_lut (.A(branch_target_d[13]), .B(bypass_data_0[13]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i12_3_lut.init = 16'hcaca;
    LUT4 mux_432_i13_3_lut (.A(branch_target_d[14]), .B(bypass_data_0[14]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i13_3_lut.init = 16'hcaca;
    LUT4 mux_432_i14_3_lut (.A(branch_target_d[15]), .B(bypass_data_0[15]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i14_3_lut.init = 16'hcaca;
    LUT4 mux_432_i15_3_lut (.A(branch_target_d[16]), .B(bypass_data_0[16]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i15_3_lut.init = 16'hcaca;
    LUT4 mux_432_i16_3_lut (.A(branch_target_d[17]), .B(bypass_data_0[17]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i16_3_lut.init = 16'hcaca;
    LUT4 mux_432_i17_3_lut (.A(branch_target_d[18]), .B(bypass_data_0[18]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i17_3_lut.init = 16'hcaca;
    LUT4 mux_432_i18_3_lut (.A(branch_target_d[19]), .B(bypass_data_0[19]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i18_3_lut.init = 16'hcaca;
    LUT4 mux_432_i19_3_lut (.A(branch_target_d[20]), .B(bypass_data_0[20]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i19_3_lut.init = 16'hcaca;
    LUT4 mux_432_i20_3_lut (.A(branch_target_d[21]), .B(bypass_data_0[21]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i20_3_lut.init = 16'hcaca;
    LUT4 mux_432_i21_3_lut (.A(branch_target_d[22]), .B(bypass_data_0[22]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i21_3_lut.init = 16'hcaca;
    LUT4 mux_432_i22_3_lut (.A(branch_target_d[23]), .B(bypass_data_0[23]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i22_3_lut.init = 16'hcaca;
    LUT4 mux_432_i23_3_lut (.A(branch_target_d[24]), .B(bypass_data_0[24]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i23_3_lut.init = 16'hcaca;
    LUT4 mux_432_i24_3_lut (.A(branch_target_d[25]), .B(bypass_data_0[25]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i24_3_lut.init = 16'hcaca;
    LUT4 mux_432_i25_3_lut (.A(branch_target_d[26]), .B(bypass_data_0[26]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i25_3_lut.init = 16'hcaca;
    LUT4 mux_432_i26_3_lut (.A(branch_target_d[27]), .B(bypass_data_0[27]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i26_3_lut.init = 16'hcaca;
    LUT4 mux_432_i27_3_lut (.A(branch_target_d[28]), .B(bypass_data_0[28]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i27_3_lut.init = 16'hcaca;
    LUT4 mux_432_i28_3_lut (.A(branch_target_d[29]), .B(bypass_data_0[29]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i28_3_lut.init = 16'hcaca;
    LUT4 mux_432_i29_3_lut (.A(branch_target_d[30]), .B(bypass_data_0[30]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i29_3_lut.init = 16'hcaca;
    LUT4 mux_432_i30_3_lut (.A(branch_target_d[31]), .B(bypass_data_0[31]), 
         .C(n6026), .Z(branch_target_x_31__N_1120[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_432_i30_3_lut.init = 16'hcaca;
    LUT4 mux_508_i4_4_lut (.A(branch_target_x[5]), .B(eid_x_2__N_1108[0]), 
         .C(n41202), .D(n41414), .Z(branch_target_m_31__N_1167[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2555[7:45])
    defparam mux_508_i4_4_lut.init = 16'h0aca;
    LUT4 i14583_4_lut (.A(n41416), .B(n41417), .C(n41415), .D(divide_by_zero_x), 
         .Z(eid_x_2__N_1108[0])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B+!(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1838[10] 1864[33])
    defparam i14583_4_lut.init = 16'hcfcd;
    LUT4 mux_508_i30_3_lut_4_lut_else_3_lut (.A(n41417), .B(deba[31]), .C(branch_target_x[31]), 
         .Z(n41498)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1795[22:86])
    defparam mux_508_i30_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 mux_508_i6_4_lut (.A(branch_target_x[7]), .B(eid_x_2__N_1009[2]), 
         .C(n41202), .D(reset_exception), .Z(branch_target_m_31__N_1167[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2555[7:45])
    defparam mux_508_i6_4_lut.init = 16'h0aca;
    LUT4 i1_2_lut_rep_1025 (.A(valid_w), .B(write_enable_w), .Z(n41430)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2700[10] 2703[12])
    defparam i1_2_lut_rep_1025.init = 16'h8888;
    LUT4 i1_3_lut_rep_920_4_lut (.A(valid_w), .B(write_enable_w), .C(\counter[2] ), 
         .D(dcache_refill_request), .Z(n41325)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2700[10] 2703[12])
    defparam i1_3_lut_rep_920_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_1088 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_442)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1088.init = 16'h0f0e;
    LUT4 condition_met_m_bdd_3_lut (.A(condition_met_m), .B(branch_predict_m), 
         .C(branch_predict_taken_m), .Z(branch_taken_m_N_1388)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;
    defparam condition_met_m_bdd_3_lut.init = 16'h4a4a;
    LUT4 i1_2_lut_rep_1124 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_456)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1124.init = 16'h0f0e;
    PFUMX i34530 (.BLUT(n41766), .ALUT(n41762), .C0(x_result_sel_csr_x), 
          .Z(n41767));
    LUT4 i1_2_lut_rep_1031 (.A(dcache_refill_request), .B(valid_m), .Z(n41436)) /* synthesis lut_function=(!(A+!(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[14:54])
    defparam i1_2_lut_rep_1031.init = 16'h4444;
    LUT4 store_m_I_0_2_lut_rep_878_3_lut_4_lut (.A(dcache_refill_request), 
         .B(valid_m), .C(store_m), .D(exception_m), .Z(n41283)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[14:54])
    defparam store_m_I_0_2_lut_rep_878_3_lut_4_lut.init = 16'h0040;
    LUT4 cmp_zero_bdd_3_lut (.A(operand_0_x[31]), .B(\adder_result_x[31] ), 
         .C(operand_1_x[31]), .Z(n40686)) /* synthesis lut_function=(!(A (B+!(C))+!A !((C)+!B))) */ ;
    defparam cmp_zero_bdd_3_lut.init = 16'h7171;
    LUT4 i1_2_lut_rep_955_3_lut (.A(dcache_refill_request), .B(valid_m), 
         .C(exception_m), .Z(n41360)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[14:54])
    defparam i1_2_lut_rep_955_3_lut.init = 16'h0404;
    LUT4 load_m_I_0_2_lut_rep_879_3_lut_4_lut (.A(dcache_refill_request), 
         .B(valid_m), .C(load_m), .D(exception_m), .Z(n41284)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[14:54])
    defparam load_m_I_0_2_lut_rep_879_3_lut_4_lut.init = 16'h0040;
    LUT4 cmp_zero_bdd_4_lut (.A(size_x[0]), .B(operand_0_x[31]), .C(\adder_result_x[31] ), 
         .D(operand_1_x[31]), .Z(n40685)) /* synthesis lut_function=(!((B (C+!(D))+!B !((D)+!C))+!A)) */ ;
    defparam cmp_zero_bdd_4_lut.init = 16'h2a02;
    LUT4 operand_w_31__I_0_i1_3_lut (.A(operand_w[0]), .B(multiplier_result_w[0]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 adder_carry_n_x_bdd_4_lut (.A(adder_carry_n_x), .B(cmp_zero), .C(size_x[0]), 
         .D(size_x[1]), .Z(n40684)) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(D)))) */ ;
    defparam adder_carry_n_x_bdd_4_lut.init = 16'h3f2a;
    LUT4 n41732_bdd_3_lut (.A(n41732), .B(adder_result_x[8]), .C(x_result_sel_add_x), 
         .Z(x_result[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41732_bdd_3_lut.init = 16'hcaca;
    LUT4 logic_result_x_9__bdd_4_lut_34507 (.A(n39318), .B(n5915), .C(n39317), 
         .D(csr_x[2]), .Z(n41734)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam logic_result_x_9__bdd_4_lut_34507.init = 16'hc088;
    LUT4 logic_result_x_9__bdd_4_lut_35823 (.A(size_x[1]), .B(size_x[0]), 
         .C(operand_0_x[9]), .D(operand_0_x[7]), .Z(n41735)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam logic_result_x_9__bdd_4_lut_35823.init = 16'hf1e0;
    LUT4 logic_result_x_9__bdd_3_lut_35824 (.A(size_x[1]), .B(size_x[0]), 
         .C(operand_0_x[9]), .Z(n41736)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam logic_result_x_9__bdd_3_lut_35824.init = 16'hacac;
    LUT4 i1_3_lut_adj_635 (.A(exception_m), .B(n41302), .C(m_result_sel_compare_m), 
         .Z(operand_w_31__N_850[1])) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i1_3_lut_adj_635.init = 16'h0404;
    LUT4 m_result_31__I_0_i3_3_lut (.A(m_result[2]), .B(operand_w_31__N_1197[2]), 
         .C(exception_m), .Z(operand_w_31__N_850[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i1_3_lut (.A(pc_m[2]), .B(memop_pc_w[2]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i1_3_lut.init = 16'hcaca;
    LUT4 i15003_4_lut (.A(operand_m[2]), .B(m_result_sel_compare_m), .C(shifter_result_m[2]), 
         .D(m_result_sel_shift_m), .Z(m_result[2])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15003_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i4_3_lut (.A(m_result[3]), .B(operand_w_31__N_1197[3]), 
         .C(exception_m), .Z(operand_w_31__N_850[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i2_3_lut (.A(pc_m[3]), .B(memop_pc_w[3]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i2_3_lut.init = 16'hcaca;
    LUT4 i15004_4_lut (.A(operand_m[3]), .B(m_result_sel_compare_m), .C(shifter_result_m[3]), 
         .D(m_result_sel_shift_m), .Z(m_result[3])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15004_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i5_3_lut (.A(m_result[4]), .B(operand_w_31__N_1197[4]), 
         .C(exception_m), .Z(operand_w_31__N_850[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i3_3_lut (.A(pc_m[4]), .B(memop_pc_w[4]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i3_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_636 (.A(m_result_sel_compare_m), .B(operand_m[4]), 
         .C(n19316), .D(m_result_sel_shift_m), .Z(m_result[4])) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i1_4_lut_adj_636.init = 16'h5044;
    LUT4 i14042_3_lut (.A(left_shift_result[27]), .B(left_shift_result[4]), 
         .C(direction_m), .Z(n19316)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(92[5:16])
    defparam i14042_3_lut.init = 16'hcaca;
    LUT4 m_result_31__I_0_i6_3_lut (.A(m_result[5]), .B(operand_w_31__N_1197[5]), 
         .C(exception_m), .Z(operand_w_31__N_850[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_1089 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_441)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1089.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_1090 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_440)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1090.init = 16'h0f0e;
    LUT4 mux_1682_i4_3_lut (.A(pc_m[5]), .B(memop_pc_w[5]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i4_3_lut.init = 16'hcaca;
    LUT4 i15005_4_lut (.A(\operand_m[5] ), .B(m_result_sel_compare_m), .C(shifter_result_m[5]), 
         .D(m_result_sel_shift_m), .Z(m_result[5])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15005_4_lut.init = 16'h3022;
    LUT4 i15416_4_lut (.A(ie), .B(n31825), .C(im[0]), .D(csr_x[0]), 
         .Z(n5814[0])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15416_4_lut.init = 16'hc088;
    LUT4 i15098_3_lut_3_lut_3_lut (.A(csr_x[3]), .B(eba[17]), .C(csr_x[0]), 
         .Z(n5780[17])) /* synthesis lut_function=(!(A+!(B+!(C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2132[5:19])
    defparam i15098_3_lut_3_lut_3_lut.init = 16'h4545;
    PFUMX i34528 (.BLUT(logic_result_x[13]), .ALUT(n41764), .C0(n36746), 
          .Z(n41765));
    LUT4 i15099_3_lut_3_lut_3_lut (.A(csr_x[3]), .B(eba[27]), .C(csr_x[0]), 
         .Z(n5780[27])) /* synthesis lut_function=(!(A+!(B+!(C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2132[5:19])
    defparam i15099_3_lut_3_lut_3_lut.init = 16'h4545;
    LUT4 n10760_bdd_2_lut_33715_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[9]), 
         .Z(n39317)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam n10760_bdd_2_lut_33715_3_lut.init = 16'h2020;
    LUT4 n10760_bdd_2_lut_33722_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[10]), 
         .Z(n39320)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam n10760_bdd_2_lut_33722_3_lut.init = 16'h2020;
    LUT4 n10760_bdd_2_lut_33744_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[14]), 
         .Z(n39332)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam n10760_bdd_2_lut_33744_3_lut.init = 16'h2020;
    LUT4 n10760_bdd_2_lut_33726_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[12]), 
         .Z(n39326)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam n10760_bdd_2_lut_33726_3_lut.init = 16'h2020;
    LUT4 n10760_bdd_2_lut_33730_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[13]), 
         .Z(n39329)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam n10760_bdd_2_lut_33730_3_lut.init = 16'h2020;
    LUT4 i15345_2_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[15]), 
         .Z(n5780[15])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15345_2_lut_3_lut.init = 16'h2020;
    LUT4 i15348_2_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[16]), 
         .Z(n5780[16])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15348_2_lut_3_lut.init = 16'h2020;
    LUT4 i15349_2_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[18]), 
         .Z(n5780[18])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15349_2_lut_3_lut.init = 16'h2020;
    LUT4 m_result_31__I_0_i7_3_lut (.A(m_result[6]), .B(operand_w_31__N_1197[6]), 
         .C(exception_m), .Z(operand_w_31__N_850[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i5_3_lut (.A(pc_m[6]), .B(memop_pc_w[6]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i5_3_lut.init = 16'hcaca;
    LUT4 i15350_2_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[19]), 
         .Z(n5780[19])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15350_2_lut_3_lut.init = 16'h2020;
    LUT4 i15351_2_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[20]), 
         .Z(n5780[20])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15351_2_lut_3_lut.init = 16'h2020;
    LUT4 i15352_2_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[21]), 
         .Z(n5780[21])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15352_2_lut_3_lut.init = 16'h2020;
    LUT4 i15353_2_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[22]), 
         .Z(n5780[22])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15353_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_4_lut_adj_637 (.A(m_result_sel_compare_m), .B(operand_m[6]), 
         .C(n19330), .D(m_result_sel_shift_m), .Z(m_result[6])) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i1_4_lut_adj_637.init = 16'h5044;
    LUT4 i14057_3_lut (.A(left_shift_result[25]), .B(left_shift_result[6]), 
         .C(direction_m), .Z(n19330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(92[5:16])
    defparam i14057_3_lut.init = 16'hcaca;
    LUT4 m_result_31__I_0_i8_3_lut (.A(m_result[7]), .B(operand_w_31__N_1197[7]), 
         .C(exception_m), .Z(operand_w_31__N_850[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 i15354_2_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[23]), 
         .Z(n5780[23])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15354_2_lut_3_lut.init = 16'h2020;
    LUT4 i15355_2_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[24]), 
         .Z(n5780[24])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15355_2_lut_3_lut.init = 16'h2020;
    LUT4 i15356_2_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[25]), 
         .Z(n5780[25])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15356_2_lut_3_lut.init = 16'h2020;
    LUT4 i15357_2_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[26]), 
         .Z(n5780[26])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15357_2_lut_3_lut.init = 16'h2020;
    LUT4 i15358_2_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[28]), 
         .Z(n5780[28])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15358_2_lut_3_lut.init = 16'h2020;
    LUT4 i15359_2_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[29]), 
         .Z(n5780[29])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15359_2_lut_3_lut.init = 16'h2020;
    LUT4 i15362_2_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[30]), 
         .Z(n5780[30])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15362_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_1091 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_439)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1091.init = 16'h0f0e;
    LUT4 i15365_2_lut_3_lut (.A(csr_x[0]), .B(csr_x[3]), .C(eba[31]), 
         .Z(n5780[31])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i15365_2_lut_3_lut.init = 16'h2020;
    LUT4 i33070_2_lut_rep_1039 (.A(x_result_sel_csr_x), .B(x_result_sel_sext_x), 
         .Z(n41444)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam i33070_2_lut_rep_1039.init = 16'heeee;
    LUT4 i1_2_lut_rep_1125 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_455)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1125.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_1126 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_454)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1126.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_1127 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_453)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1127.init = 16'h0f0e;
    LUT4 mux_1682_i6_3_lut (.A(pc_m[7]), .B(memop_pc_w[7]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i6_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_1128 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_452)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1128.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_1129 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_451)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1129.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_1130 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_450)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1130.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_1131 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_449)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1131.init = 16'h0f0e;
    LUT4 i15006_4_lut (.A(operand_m[7]), .B(m_result_sel_compare_m), .C(shifter_result_m[7]), 
         .D(m_result_sel_shift_m), .Z(m_result[7])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15006_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i9_3_lut (.A(m_result[8]), .B(operand_w_31__N_1197[8]), 
         .C(exception_m), .Z(operand_w_31__N_850[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 n10760_bdd_4_lut_33719 (.A(n41288), .B(n41391), .C(im[10]), .D(deba[10]), 
         .Z(n39321)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (D))) */ ;
    defparam n10760_bdd_4_lut_33719.init = 16'hec20;
    LUT4 mux_1682_i7_3_lut (.A(pc_m[8]), .B(memop_pc_w[8]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i7_3_lut.init = 16'hcaca;
    LUT4 i15007_4_lut (.A(operand_m[8]), .B(m_result_sel_compare_m), .C(shifter_result_m[8]), 
         .D(m_result_sel_shift_m), .Z(m_result[8])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15007_4_lut.init = 16'h3022;
    LUT4 i15108_2_lut_2_lut (.A(dcache_refill_request), .B(operand_m[2]), 
         .Z(d_adr_o_31__N_2278[2])) /* synthesis lut_function=(!(A+!(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[36:54])
    defparam i15108_2_lut_2_lut.init = 16'h4444;
    LUT4 i15109_2_lut_2_lut (.A(dcache_refill_request), .B(operand_m[3]), 
         .Z(d_adr_o_31__N_2278[3])) /* synthesis lut_function=(!(A+!(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[36:54])
    defparam i15109_2_lut_2_lut.init = 16'h4444;
    LUT4 m_result_31__I_0_i10_3_lut (.A(m_result[9]), .B(operand_w_31__N_1197[9]), 
         .C(exception_m), .Z(operand_w_31__N_850[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i8_3_lut (.A(pc_m[9]), .B(memop_pc_w[9]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i8_3_lut.init = 16'hcaca;
    LUT4 i15008_4_lut (.A(\operand_m[9] ), .B(m_result_sel_compare_m), .C(shifter_result_m[9]), 
         .D(m_result_sel_shift_m), .Z(m_result[9])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15008_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i11_3_lut (.A(m_result[10]), .B(operand_w_31__N_1197[10]), 
         .C(exception_m), .Z(operand_w_31__N_850[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i9_3_lut (.A(pc_m[10]), .B(memop_pc_w[10]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i9_3_lut.init = 16'hcaca;
    LUT4 i15009_4_lut (.A(\operand_m[10] ), .B(m_result_sel_compare_m), 
         .C(n17816), .D(m_result_sel_shift_m), .Z(m_result[10])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15009_4_lut.init = 16'h3022;
    LUT4 i30443_2_lut_3_lut_4_lut (.A(write_idx_m[2]), .B(n41359), .C(n41358), 
         .D(write_idx_m[1]), .Z(n35587)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1489[18:47])
    defparam i30443_2_lut_3_lut_4_lut.init = 16'h6ff6;
    LUT4 m_result_31__I_0_i12_3_lut (.A(m_result[11]), .B(operand_w_31__N_1197[11]), 
         .C(exception_m), .Z(operand_w_31__N_850[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i10_3_lut (.A(pc_m[11]), .B(memop_pc_w[11]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i10_3_lut.init = 16'hcaca;
    LUT4 i15010_4_lut (.A(operand_m[11]), .B(m_result_sel_compare_m), .C(shifter_result_m[11]), 
         .D(m_result_sel_shift_m), .Z(m_result[11])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15010_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i13_3_lut (.A(m_result[12]), .B(operand_w_31__N_1197[12]), 
         .C(exception_m), .Z(operand_w_31__N_850[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i11_3_lut (.A(pc_m[12]), .B(memop_pc_w[12]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i11_3_lut.init = 16'hcaca;
    LUT4 i14688_2_lut_3_lut_4_lut (.A(store_m), .B(n41360), .C(n41389), 
         .D(n45171), .Z(n12404)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2005[20:56])
    defparam i14688_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_638 (.A(store_m), .B(n41360), .C(n20639), 
         .D(n45171), .Z(REF_CLK_c_enable_949)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2005[20:56])
    defparam i1_2_lut_3_lut_4_lut_adj_638.init = 16'h0800;
    LUT4 i15011_4_lut (.A(operand_m[12]), .B(m_result_sel_compare_m), .C(shifter_result_m[12]), 
         .D(m_result_sel_shift_m), .Z(m_result[12])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15011_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i14_3_lut (.A(m_result[13]), .B(operand_w_31__N_1197[13]), 
         .C(exception_m), .Z(operand_w_31__N_850[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i12_3_lut (.A(pc_m[13]), .B(memop_pc_w[13]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i12_3_lut.init = 16'hcaca;
    LUT4 i15012_4_lut (.A(operand_m[13]), .B(m_result_sel_compare_m), .C(shifter_result_m[13]), 
         .D(m_result_sel_shift_m), .Z(m_result[13])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15012_4_lut.init = 16'h3022;
    LUT4 csr_x_4__I_0_738_i7_2_lut_rep_1043 (.A(csr_x[3]), .B(csr_x[4]), 
         .Z(n41448)) /* synthesis lut_function=((B)+!A) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2132[5:19])
    defparam csr_x_4__I_0_738_i7_2_lut_rep_1043.init = 16'hdddd;
    LUT4 m_result_31__I_0_i15_3_lut (.A(m_result[14]), .B(operand_w_31__N_1197[14]), 
         .C(exception_m), .Z(operand_w_31__N_850[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i15_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_639 (.A(csr_x[3]), .B(csr_x[4]), .C(n41449), 
         .D(csr_x[2]), .Z(n34890)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2132[5:19])
    defparam i1_2_lut_3_lut_4_lut_adj_639.init = 16'h0020;
    LUT4 mux_1682_i13_3_lut (.A(pc_m[14]), .B(memop_pc_w[14]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i13_3_lut.init = 16'hcaca;
    PFUMX i34353 (.BLUT(n41166), .ALUT(n41165), .C0(w_result_sel_load_w), 
          .Z(w_result[8]));
    LUT4 i15319_2_lut_rep_974_3_lut (.A(csr_x[3]), .B(csr_x[4]), .C(csr_x[2]), 
         .Z(n41379)) /* synthesis lut_function=((B+(C))+!A) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2132[5:19])
    defparam i15319_2_lut_rep_974_3_lut.init = 16'hfdfd;
    LUT4 i1_2_lut_rep_1044 (.A(csr_x[1]), .B(csr_x[0]), .Z(n41449)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_rep_1044.init = 16'h4444;
    LUT4 i15013_4_lut (.A(operand_m[14]), .B(m_result_sel_compare_m), .C(shifter_result_m[14]), 
         .D(m_result_sel_shift_m), .Z(m_result[14])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15013_4_lut.init = 16'h3022;
    LUT4 i1_3_lut_4_lut_adj_640 (.A(store_m), .B(n41360), .C(dcache_select_m), 
         .D(state_adj_6256[1]), .Z(n30107)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2005[20:56])
    defparam i1_3_lut_4_lut_adj_640.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_641 (.A(csr_x[1]), .B(csr_x[0]), .C(valid_w), 
         .D(debug_exception_w), .Z(n34874)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_641.init = 16'h0444;
    LUT4 i1_2_lut_rep_1045 (.A(branch_predict_taken_m), .B(branch_predict_m), 
         .Z(n41450)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i1_2_lut_rep_1045.init = 16'h8888;
    LUT4 i1_2_lut_rep_944_3_lut (.A(branch_predict_taken_m), .B(branch_predict_m), 
         .C(condition_met_m), .Z(n41349)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i1_2_lut_rep_944_3_lut.init = 16'h0808;
    LUT4 m_result_31__I_0_i16_3_lut (.A(m_result[15]), .B(operand_w_31__N_1197[15]), 
         .C(exception_m), .Z(operand_w_31__N_850[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i16_3_lut.init = 16'hcaca;
    LUT4 n10760_bdd_4_lut_33716 (.A(n41288), .B(n41391), .C(im[9]), .D(deba[9]), 
         .Z(n39318)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (D))) */ ;
    defparam n10760_bdd_4_lut_33716.init = 16'hec20;
    LUT4 i1_3_lut_rep_810_4_lut (.A(load_m), .B(n41360), .C(wb_select_m), 
         .D(wb_load_complete), .Z(n41215)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2004[19:54])
    defparam i1_3_lut_rep_810_4_lut.init = 16'h0080;
    LUT4 mux_1682_i14_3_lut (.A(pc_m[15]), .B(memop_pc_w[15]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i14_3_lut.init = 16'hcaca;
    LUT4 i15014_4_lut (.A(operand_m[15]), .B(m_result_sel_compare_m), .C(shifter_result_m[15]), 
         .D(m_result_sel_shift_m), .Z(m_result[15])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15014_4_lut.init = 16'h3022;
    LUT4 i1_3_lut_4_lut_4_lut (.A(load_m), .B(n41360), .C(LM32D_CYC_O), 
         .D(store_m), .Z(n32408)) /* synthesis lut_function=(A (B+(C))+!A (B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2004[19:54])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hfcf8;
    PFUMX i34525 (.BLUT(n41759), .ALUT(n41755), .C0(x_result_sel_csr_x), 
          .Z(n41760));
    LUT4 m_result_31__I_0_i17_3_lut (.A(m_result[16]), .B(operand_w_31__N_1197[16]), 
         .C(exception_m), .Z(operand_w_31__N_850[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i15_3_lut (.A(pc_m[16]), .B(memop_pc_w[16]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i15_3_lut.init = 16'hcaca;
    LUT4 i15015_4_lut (.A(operand_m[16]), .B(m_result_sel_compare_m), .C(shifter_result_m[16]), 
         .D(m_result_sel_shift_m), .Z(m_result[16])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15015_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i18_3_lut (.A(m_result[17]), .B(operand_w_31__N_1197[17]), 
         .C(exception_m), .Z(operand_w_31__N_850[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i16_3_lut (.A(pc_m[17]), .B(memop_pc_w[17]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i16_3_lut.init = 16'hcaca;
    LUT4 i15016_4_lut (.A(operand_m[17]), .B(m_result_sel_compare_m), .C(shifter_result_m[17]), 
         .D(m_result_sel_shift_m), .Z(m_result[17])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15016_4_lut.init = 16'h3022;
    PFUMX i34523 (.BLUT(logic_result_x[12]), .ALUT(n41757), .C0(n36735), 
          .Z(n41758));
    LUT4 m_result_31__I_0_i19_3_lut (.A(m_result[18]), .B(operand_w_31__N_1197[18]), 
         .C(exception_m), .Z(operand_w_31__N_850[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i19_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i17_3_lut (.A(pc_m[18]), .B(memop_pc_w[18]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i17_3_lut.init = 16'hcaca;
    PFUMX i34520 (.BLUT(n41752), .ALUT(n41748), .C0(x_result_sel_csr_x), 
          .Z(n41753));
    PFUMX i34348 (.BLUT(n41162), .ALUT(n41161), .C0(w_result_sel_load_w), 
          .Z(w_result[9]));
    LUT4 i15017_4_lut (.A(operand_m[18]), .B(m_result_sel_compare_m), .C(shifter_result_m[18]), 
         .D(m_result_sel_shift_m), .Z(m_result[18])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15017_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i20_3_lut (.A(m_result[19]), .B(operand_w_31__N_1197[19]), 
         .C(exception_m), .Z(operand_w_31__N_850[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i18_3_lut (.A(pc_m[19]), .B(memop_pc_w[19]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i18_3_lut.init = 16'hcaca;
    LUT4 i15018_4_lut (.A(operand_m[19]), .B(m_result_sel_compare_m), .C(shifter_result_m[19]), 
         .D(m_result_sel_shift_m), .Z(m_result[19])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15018_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i21_3_lut (.A(m_result[20]), .B(operand_w_31__N_1197[20]), 
         .C(exception_m), .Z(operand_w_31__N_850[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i19_3_lut (.A(pc_m[20]), .B(memop_pc_w[20]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i19_3_lut.init = 16'hcaca;
    LUT4 i15019_4_lut (.A(operand_m[20]), .B(m_result_sel_compare_m), .C(shifter_result_m[20]), 
         .D(m_result_sel_shift_m), .Z(m_result[20])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15019_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i22_3_lut (.A(m_result[21]), .B(operand_w_31__N_1197[21]), 
         .C(exception_m), .Z(operand_w_31__N_850[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i22_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i20_3_lut (.A(pc_m[21]), .B(memop_pc_w[21]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i20_3_lut.init = 16'hcaca;
    LUT4 i15020_4_lut (.A(operand_m[21]), .B(m_result_sel_compare_m), .C(\shifter_result_m[21] ), 
         .D(m_result_sel_shift_m), .Z(m_result[21])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15020_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i23_3_lut (.A(m_result[22]), .B(operand_w_31__N_1197[22]), 
         .C(exception_m), .Z(operand_w_31__N_850[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i23_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i21_3_lut (.A(pc_m[22]), .B(memop_pc_w[22]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i21_3_lut.init = 16'hcaca;
    LUT4 i15021_4_lut (.A(operand_m[22]), .B(m_result_sel_compare_m), .C(shifter_result_m[22]), 
         .D(m_result_sel_shift_m), .Z(m_result[22])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15021_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i24_3_lut (.A(m_result[23]), .B(operand_w_31__N_1197[23]), 
         .C(exception_m), .Z(operand_w_31__N_850[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i24_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i22_3_lut (.A(pc_m[23]), .B(memop_pc_w[23]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i22_3_lut.init = 16'hcaca;
    LUT4 i15022_4_lut (.A(operand_m[23]), .B(m_result_sel_compare_m), .C(shifter_result_m[23]), 
         .D(m_result_sel_shift_m), .Z(m_result[23])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15022_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i25_3_lut (.A(m_result[24]), .B(operand_w_31__N_1197[24]), 
         .C(exception_m), .Z(operand_w_31__N_850[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i25_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i23_3_lut (.A(pc_m[24]), .B(memop_pc_w[24]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i23_3_lut.init = 16'hcaca;
    LUT4 i15023_4_lut (.A(operand_m[24]), .B(m_result_sel_compare_m), .C(shifter_result_m[24]), 
         .D(m_result_sel_shift_m), .Z(m_result[24])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15023_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i26_3_lut (.A(m_result[25]), .B(operand_w_31__N_1197[25]), 
         .C(exception_m), .Z(operand_w_31__N_850[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i26_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i24_3_lut (.A(pc_m[25]), .B(memop_pc_w[25]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i24_3_lut.init = 16'hcaca;
    LUT4 i15024_4_lut (.A(operand_m[25]), .B(m_result_sel_compare_m), .C(n19333), 
         .D(m_result_sel_shift_m), .Z(m_result[25])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15024_4_lut.init = 16'h3022;
    LUT4 i14060_3_lut (.A(left_shift_result[6]), .B(left_shift_result[25]), 
         .C(direction_m), .Z(n19333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(92[5:16])
    defparam i14060_3_lut.init = 16'hcaca;
    LUT4 m_result_31__I_0_i27_3_lut (.A(m_result[26]), .B(operand_w_31__N_1197[26]), 
         .C(exception_m), .Z(operand_w_31__N_850[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i27_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i25_3_lut (.A(pc_m[26]), .B(memop_pc_w[26]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i25_3_lut.init = 16'hcaca;
    LUT4 i15025_4_lut (.A(operand_m[26]), .B(m_result_sel_compare_m), .C(shifter_result_m[26]), 
         .D(m_result_sel_shift_m), .Z(m_result[26])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15025_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i28_3_lut (.A(m_result[27]), .B(operand_w_31__N_1197[27]), 
         .C(exception_m), .Z(operand_w_31__N_850[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i28_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i26_3_lut (.A(pc_m[27]), .B(memop_pc_w[27]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i26_3_lut.init = 16'hcaca;
    LUT4 i15026_4_lut (.A(operand_m[27]), .B(m_result_sel_compare_m), .C(n19319), 
         .D(m_result_sel_shift_m), .Z(m_result[27])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15026_4_lut.init = 16'h3022;
    LUT4 i14045_3_lut (.A(left_shift_result[4]), .B(left_shift_result[27]), 
         .C(direction_m), .Z(n19319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(92[5:16])
    defparam i14045_3_lut.init = 16'hcaca;
    LUT4 m_result_31__I_0_i29_3_lut (.A(m_result[28]), .B(operand_w_31__N_1197[28]), 
         .C(exception_m), .Z(operand_w_31__N_850[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i29_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i27_3_lut (.A(pc_m[28]), .B(memop_pc_w[28]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i27_3_lut.init = 16'hcaca;
    LUT4 i15027_4_lut (.A(operand_m[28]), .B(m_result_sel_compare_m), .C(shifter_result_m[28]), 
         .D(m_result_sel_shift_m), .Z(m_result[28])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15027_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i30_3_lut (.A(m_result[29]), .B(operand_w_31__N_1197[29]), 
         .C(exception_m), .Z(operand_w_31__N_850[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i30_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i28_3_lut (.A(pc_m[29]), .B(memop_pc_w[29]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i28_3_lut.init = 16'hcaca;
    LUT4 i15028_4_lut (.A(operand_m[29]), .B(m_result_sel_compare_m), .C(shifter_result_m[29]), 
         .D(m_result_sel_shift_m), .Z(m_result[29])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15028_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i31_3_lut (.A(m_result[30]), .B(operand_w_31__N_1197[30]), 
         .C(exception_m), .Z(operand_w_31__N_850[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i31_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i29_3_lut (.A(pc_m[30]), .B(memop_pc_w[30]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i29_3_lut.init = 16'hcaca;
    PFUMX i34343 (.BLUT(n41158), .ALUT(n41157), .C0(w_result_sel_load_w), 
          .Z(w_result[10]));
    LUT4 i15029_4_lut (.A(operand_m[30]), .B(m_result_sel_compare_m), .C(shifter_result_m[30]), 
         .D(m_result_sel_shift_m), .Z(m_result[30])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15029_4_lut.init = 16'h3022;
    LUT4 m_result_31__I_0_i32_3_lut (.A(m_result[31]), .B(operand_w_31__N_1197[31]), 
         .C(exception_m), .Z(operand_w_31__N_850[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i32_3_lut.init = 16'hcaca;
    LUT4 mux_1682_i30_3_lut (.A(pc_m[31]), .B(memop_pc_w[31]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1197[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_1682_i30_3_lut.init = 16'hcaca;
    LUT4 i15030_4_lut (.A(operand_m[31]), .B(m_result_sel_compare_m), .C(shifter_result_m[31]), 
         .D(m_result_sel_shift_m), .Z(m_result[31])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i15030_4_lut.init = 16'h3022;
    LUT4 i12666_3_lut (.A(left_shift_result[0]), .B(left_shift_result[31]), 
         .C(direction_m), .Z(shifter_result_m[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(92[5:16])
    defparam i12666_3_lut.init = 16'hcaca;
    PFUMX i34338 (.BLUT(n41154), .ALUT(n41153), .C0(w_result_sel_load_w), 
          .Z(w_result[11]));
    LUT4 logic_result_x_8__bdd_3_lut_34552 (.A(size_x[1]), .B(size_x[0]), 
         .C(operand_0_x[8]), .Z(n41729)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam logic_result_x_8__bdd_3_lut_34552.init = 16'hacac;
    LUT4 bypass_data_0_31__I_14_i2_3_lut_4_lut (.A(n41302), .B(m_result_sel_compare_m), 
         .C(raw_x_0), .D(x_result[1]), .Z(bypass_data_0_31__N_882[1])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam bypass_data_0_31__I_14_i2_3_lut_4_lut.init = 16'hf202;
    LUT4 bypass_data_1_31__I_15_i2_3_lut_4_lut (.A(n41302), .B(m_result_sel_compare_m), 
         .C(raw_x_1), .D(x_result[1]), .Z(bypass_data_1_31__N_914[1])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam bypass_data_1_31__I_15_i2_3_lut_4_lut.init = 16'hf202;
    PFUMX i34333 (.BLUT(n41150), .ALUT(n41149), .C0(w_result_sel_load_w), 
          .Z(w_result[12]));
    PFUMX i34328 (.BLUT(n41146), .ALUT(n41145), .C0(w_result_sel_load_w), 
          .Z(w_result[13]));
    LUT4 eba_8__bdd_3_lut (.A(\jtag_reg_addr_d[0] ), .B(\jtag_reg_addr_d[1] ), 
         .C(csr_x[0]), .Z(n39310)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam eba_8__bdd_3_lut.init = 16'hcaca;
    LUT4 mux_13_i26_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[27]), 
         .D(branch_target_m[27]), .Z(pc_a_31__N_1720[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i26_3_lut_4_lut.init = 16'hfd20;
    LUT4 n40688_bdd_3_lut_4_lut (.A(cmp_zero), .B(size_x[0]), .C(size_x[1]), 
         .D(n40687), .Z(n40689)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam n40688_bdd_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_13_i27_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[28]), 
         .D(branch_target_m[28]), .Z(pc_a_31__N_1720[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i27_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i28_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[29]), 
         .D(branch_target_m[29]), .Z(pc_a_31__N_1720[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i28_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i29_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[30]), 
         .D(branch_target_m[30]), .Z(pc_a_31__N_1720[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i29_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i30_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[31]), 
         .D(branch_target_m[31]), .Z(pc_a_31__N_1720[29])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i30_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i7_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[8]), 
         .D(branch_target_m[8]), .Z(pc_a_31__N_1720[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i5_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[6]), 
         .D(branch_target_m[6]), .Z(pc_a_31__N_1720[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_rep_1092 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_438)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1092.init = 16'h0f0e;
    LUT4 mux_13_i3_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[4]), 
         .D(branch_target_m[4]), .Z(pc_a_31__N_1720[2])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i3_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i6_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[7]), 
         .D(branch_target_m[7]), .Z(pc_a_31__N_1720[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i8_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[9]), 
         .D(branch_target_m[9]), .Z(pc_a_31__N_1720[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i8_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i25_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[26]), 
         .D(branch_target_m[26]), .Z(pc_a_31__N_1720[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i25_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i24_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[25]), 
         .D(branch_target_m[25]), .Z(pc_a_31__N_1720[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i24_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i23_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[24]), 
         .D(branch_target_m[24]), .Z(pc_a_31__N_1720[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i23_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i22_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[23]), 
         .D(branch_target_m[23]), .Z(pc_a_31__N_1720[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i22_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i21_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[22]), 
         .D(branch_target_m[22]), .Z(pc_a_31__N_1720[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i21_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i20_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[21]), 
         .D(branch_target_m[21]), .Z(pc_a_31__N_1720[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i20_3_lut_4_lut.init = 16'hfd20;
    PFUMX i34323 (.BLUT(n41142), .ALUT(n41141), .C0(w_result_sel_load_w), 
          .Z(w_result[14]));
    LUT4 mux_13_i19_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[20]), 
         .D(branch_target_m[20]), .Z(pc_a_31__N_1720[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i19_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i18_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[19]), 
         .D(branch_target_m[19]), .Z(pc_a_31__N_1720[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i18_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i17_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[18]), 
         .D(branch_target_m[18]), .Z(pc_a_31__N_1720[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i16_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[17]), 
         .D(branch_target_m[17]), .Z(pc_a_31__N_1720[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i16_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i15_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[16]), 
         .D(branch_target_m[16]), .Z(pc_a_31__N_1720[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i14_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[15]), 
         .D(branch_target_m[15]), .Z(pc_a_31__N_1720[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i13_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[14]), 
         .D(branch_target_m[14]), .Z(pc_a_31__N_1720[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i12_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[13]), 
         .D(branch_target_m[13]), .Z(pc_a_31__N_1720[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i11_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[12]), 
         .D(branch_target_m[12]), .Z(pc_a_31__N_1720[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i11_3_lut_4_lut.init = 16'hfd20;
    PFUMX d_result_sel_1_d_1__I_0_Mux_25_i3 (.BLUT(n31307), .ALUT(n2_adj_6206), 
          .C0(n37939), .Z(d_result_1[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_26_i3 (.BLUT(n31305), .ALUT(n2_adj_6205), 
          .C0(n37939), .Z(d_result_1[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_27_i3 (.BLUT(n31303), .ALUT(n2_adj_6216), 
          .C0(n37939), .Z(d_result_1[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_28_i3 (.BLUT(n31301), .ALUT(n2_adj_6217), 
          .C0(d_result_sel_1_d[1]), .Z(d_result_1[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_29_i3 (.BLUT(n31299), .ALUT(n2_adj_6218), 
          .C0(d_result_sel_1_d[1]), .Z(d_result_1[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_30_i3 (.BLUT(n31297), .ALUT(n2_adj_6219), 
          .C0(d_result_sel_1_d[1]), .Z(d_result_1[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_31_i3 (.BLUT(n31324), .ALUT(n31335), 
          .C0(d_result_sel_1_d[1]), .Z(d_result_1[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_13_i10_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[11]), 
         .D(branch_target_m[11]), .Z(pc_a_31__N_1720[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i9_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[10]), 
         .D(branch_target_m[10]), .Z(pc_a_31__N_1720[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i9_3_lut_4_lut.init = 16'hfd20;
    PFUMX d_result_sel_1_d_1__I_0_Mux_1_i3 (.BLUT(n31312), .ALUT(n31215), 
          .C0(n37933), .Z(d_result_1[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_2_lut_rep_1093 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_437)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1093.init = 16'h0f0e;
    PFUMX d_result_sel_1_d_1__I_0_Mux_3_i3 (.BLUT(n31325), .ALUT(n31210), 
          .C0(n37933), .Z(d_result_1[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_13_i4_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[5]), 
         .D(branch_target_m[5]), .Z(pc_a_31__N_1720[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i4_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_13_i2_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[3]), 
         .D(branch_target_m[3]), .Z(pc_a_31__N_1720[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i2_3_lut_4_lut.init = 16'hfd20;
    PFUMX d_result_sel_1_d_1__I_0_Mux_4_i3 (.BLUT(n31294), .ALUT(n31211), 
          .C0(n37934), .Z(d_result_1[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_13_i1_3_lut_4_lut (.A(n41349), .B(exception_m), .C(pc_x[2]), 
         .D(branch_target_m[2]), .Z(pc_a_31__N_1720[0])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam mux_13_i1_3_lut_4_lut.init = 16'hfd20;
    PFUMX d_result_sel_1_d_1__I_0_Mux_5_i3 (.BLUT(n31308), .ALUT(n31209), 
          .C0(n37934), .Z(d_result_1[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_2_lut_rep_1094 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_436)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1094.init = 16'h0f0e;
    PFUMX d_result_sel_1_d_1__I_0_Mux_6_i3 (.BLUT(n31318), .ALUT(n31207), 
          .C0(n37934), .Z(d_result_1[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_7_i3 (.BLUT(n31314), .ALUT(n31214), 
          .C0(n37934), .Z(d_result_1[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_15_i3 (.BLUT(n31296), .ALUT(n31206), 
          .C0(n37936), .Z(d_result_1[15])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_16_i3 (.BLUT(n31321), .ALUT(n2_adj_6204), 
          .C0(n37937), .Z(d_result_1[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_17_i3 (.BLUT(n31319), .ALUT(n2_adj_6203), 
          .C0(n37937), .Z(d_result_1[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_18_i3 (.BLUT(n31315), .ALUT(n2_adj_6202), 
          .C0(n37937), .Z(d_result_1[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_19_i3 (.BLUT(n31313), .ALUT(n2_adj_6201), 
          .C0(n37937), .Z(d_result_1[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_20_i3 (.BLUT(n31311), .ALUT(n2_adj_6200), 
          .C0(n37938), .Z(d_result_1[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_21_i3 (.BLUT(n31295), .ALUT(n2_adj_6199), 
          .C0(n37938), .Z(d_result_1[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_22_i3 (.BLUT(n31306), .ALUT(n2_adj_6198), 
          .C0(n37938), .Z(d_result_1[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_23_i3 (.BLUT(n31317), .ALUT(n2_adj_6197), 
          .C0(n37938), .Z(d_result_1[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_24_i3 (.BLUT(n31320), .ALUT(n2_adj_6196), 
          .C0(n37939), .Z(d_result_1[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_2_lut_rep_1132 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_448)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1132.init = 16'h0f0e;
    LUT4 n10760_bdd_4_lut_33723 (.A(n41288), .B(n41391), .C(im[11]), .D(deba[11]), 
         .Z(n39324)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (D))) */ ;
    defparam n10760_bdd_4_lut_33723.init = 16'hec20;
    LUT4 i1_2_lut_rep_1133 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_447)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1133.init = 16'h0f0e;
    PFUMX d_result_sel_1_d_1__I_0_Mux_0_i3 (.BLUT(n31309), .ALUT(n31217), 
          .C0(n37933), .Z(d_result_1[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_2_i3 (.BLUT(n31310), .ALUT(n31213), 
          .C0(n37933), .Z(d_result_1[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_8_i3 (.BLUT(n31304), .ALUT(n31220), 
          .C0(n37935), .Z(d_result_1[8])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_9_i3 (.BLUT(n31316), .ALUT(n31212), 
          .C0(n37935), .Z(d_result_1[9])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_10_i3 (.BLUT(n31302), .ALUT(n31216), 
          .C0(n37935), .Z(d_result_1[10])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_11_i3 (.BLUT(n31322), .ALUT(n31221), 
          .C0(n37935), .Z(d_result_1[11])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i33277_2_lut (.A(m_result_sel_compare_m), .B(m_result_sel_shift_m), 
         .Z(n37174)) /* synthesis lut_function=(A+!(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(439[5:27])
    defparam i33277_2_lut.init = 16'hbbbb;
    PFUMX d_result_sel_1_d_1__I_0_Mux_12_i3 (.BLUT(n31300), .ALUT(n31219), 
          .C0(n37936), .Z(d_result_1[12])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_13_i3 (.BLUT(n31298), .ALUT(n31218), 
          .C0(n37936), .Z(d_result_1[13])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX d_result_sel_1_d_1__I_0_Mux_14_i3 (.BLUT(n31323), .ALUT(n31208), 
          .C0(n37936), .Z(d_result_1[14])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX i34318 (.BLUT(n41138), .ALUT(n41137), .C0(w_result_sel_load_w), 
          .Z(w_result[15]));
    PFUMX bypass_data_1_31__I_0_i32 (.BLUT(bypass_data_1_31__N_1044[31]), 
          .ALUT(bypass_data_1_31__N_914[31]), .C0(n37940), .Z(bypass_data_1[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i31 (.BLUT(bypass_data_1_31__N_1044[30]), 
          .ALUT(bypass_data_1_31__N_914[30]), .C0(n37944), .Z(bypass_data_1[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i30 (.BLUT(bypass_data_1_31__N_1044[29]), 
          .ALUT(bypass_data_1_31__N_914[29]), .C0(n37946), .Z(bypass_data_1[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i29 (.BLUT(bypass_data_1_31__N_1044[28]), 
          .ALUT(bypass_data_1_31__N_914[28]), .C0(n37942), .Z(bypass_data_1[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i28 (.BLUT(bypass_data_1_31__N_1044[27]), 
          .ALUT(bypass_data_1_31__N_914[27]), .C0(n37943), .Z(bypass_data_1[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i27 (.BLUT(bypass_data_1_31__N_1044[26]), 
          .ALUT(bypass_data_1_31__N_914[26]), .C0(n36614), .Z(bypass_data_1[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i26 (.BLUT(bypass_data_1_31__N_1044[25]), 
          .ALUT(bypass_data_1_31__N_914[25]), .C0(n37945), .Z(bypass_data_1[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i25 (.BLUT(bypass_data_1_31__N_1044[24]), 
          .ALUT(bypass_data_1_31__N_914[24]), .C0(n37941), .Z(bypass_data_1[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i24 (.BLUT(bypass_data_1_31__N_1044[23]), 
          .ALUT(bypass_data_1_31__N_914[23]), .C0(n37941), .Z(bypass_data_1[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i23 (.BLUT(bypass_data_1_31__N_1044[22]), 
          .ALUT(bypass_data_1_31__N_914[22]), .C0(n37945), .Z(bypass_data_1[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i22 (.BLUT(bypass_data_1_31__N_1044[21]), 
          .ALUT(bypass_data_1_31__N_914[21]), .C0(n36614), .Z(bypass_data_1[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i21 (.BLUT(bypass_data_1_31__N_1044[20]), 
          .ALUT(bypass_data_1_31__N_914[20]), .C0(n37943), .Z(bypass_data_1[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i20 (.BLUT(bypass_data_1_31__N_1044[19]), 
          .ALUT(bypass_data_1_31__N_914[19]), .C0(n37942), .Z(bypass_data_1[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i19 (.BLUT(bypass_data_1_31__N_1044[18]), 
          .ALUT(bypass_data_1_31__N_914[18]), .C0(n37946), .Z(bypass_data_1[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i18 (.BLUT(bypass_data_1_31__N_1044[17]), 
          .ALUT(bypass_data_1_31__N_914[17]), .C0(n37944), .Z(bypass_data_1[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i17 (.BLUT(bypass_data_1_31__N_1044[16]), 
          .ALUT(bypass_data_1_31__N_914[16]), .C0(n37940), .Z(bypass_data_1[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i16 (.BLUT(bypass_data_1_31__N_1044[15]), 
          .ALUT(bypass_data_1_31__N_914[15]), .C0(n37940), .Z(bypass_data_1[15])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i8 (.BLUT(bypass_data_1_31__N_1044[7]), .ALUT(bypass_data_1_31__N_914[7]), 
          .C0(n37941), .Z(bypass_data_1[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i7 (.BLUT(bypass_data_1_31__N_1044[6]), .ALUT(bypass_data_1_31__N_914[6]), 
          .C0(n37945), .Z(bypass_data_1[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i6 (.BLUT(bypass_data_1_31__N_1044[5]), .ALUT(bypass_data_1_31__N_914[5]), 
          .C0(n36614), .Z(bypass_data_1[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i5 (.BLUT(bypass_data_1_31__N_1044[4]), .ALUT(bypass_data_1_31__N_914[4]), 
          .C0(n37943), .Z(bypass_data_1[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i4 (.BLUT(bypass_data_1_31__N_1044[3]), .ALUT(bypass_data_1_31__N_914[3]), 
          .C0(n37942), .Z(bypass_data_1[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i3 (.BLUT(bypass_data_1_31__N_1044[2]), .ALUT(bypass_data_1_31__N_914[2]), 
          .C0(n37946), .Z(bypass_data_1[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i2 (.BLUT(bypass_data_1_31__N_1044[1]), .ALUT(bypass_data_1_31__N_914[1]), 
          .C0(n37944), .Z(bypass_data_1[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i32 (.BLUT(bypass_data_0_31__N_1012[31]), 
          .ALUT(bypass_data_0_31__N_882[31]), .C0(n37947), .Z(bypass_data_0[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i31 (.BLUT(bypass_data_0_31__N_1012[30]), 
          .ALUT(bypass_data_0_31__N_882[30]), .C0(n37951), .Z(bypass_data_0[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i30 (.BLUT(bypass_data_0_31__N_1012[29]), 
          .ALUT(bypass_data_0_31__N_882[29]), .C0(n37953), .Z(bypass_data_0[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i29 (.BLUT(bypass_data_0_31__N_1012[28]), 
          .ALUT(bypass_data_0_31__N_882[28]), .C0(n37949), .Z(bypass_data_0[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i28 (.BLUT(bypass_data_0_31__N_1012[27]), 
          .ALUT(bypass_data_0_31__N_882[27]), .C0(n37950), .Z(bypass_data_0[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i27 (.BLUT(bypass_data_0_31__N_1012[26]), 
          .ALUT(bypass_data_0_31__N_882[26]), .C0(n36552), .Z(bypass_data_0[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i26 (.BLUT(bypass_data_0_31__N_1012[25]), 
          .ALUT(bypass_data_0_31__N_882[25]), .C0(n37952), .Z(bypass_data_0[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i25 (.BLUT(bypass_data_0_31__N_1012[24]), 
          .ALUT(bypass_data_0_31__N_882[24]), .C0(n37948), .Z(bypass_data_0[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i24 (.BLUT(bypass_data_0_31__N_1012[23]), 
          .ALUT(bypass_data_0_31__N_882[23]), .C0(n37948), .Z(bypass_data_0[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i23 (.BLUT(bypass_data_0_31__N_1012[22]), 
          .ALUT(bypass_data_0_31__N_882[22]), .C0(n37952), .Z(bypass_data_0[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i22 (.BLUT(bypass_data_0_31__N_1012[21]), 
          .ALUT(bypass_data_0_31__N_882[21]), .C0(n36552), .Z(bypass_data_0[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i21 (.BLUT(bypass_data_0_31__N_1012[20]), 
          .ALUT(bypass_data_0_31__N_882[20]), .C0(n37950), .Z(bypass_data_0[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i20 (.BLUT(bypass_data_0_31__N_1012[19]), 
          .ALUT(bypass_data_0_31__N_882[19]), .C0(n37949), .Z(bypass_data_0[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i19 (.BLUT(bypass_data_0_31__N_1012[18]), 
          .ALUT(bypass_data_0_31__N_882[18]), .C0(n37953), .Z(bypass_data_0[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i18 (.BLUT(bypass_data_0_31__N_1012[17]), 
          .ALUT(bypass_data_0_31__N_882[17]), .C0(n37951), .Z(bypass_data_0[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i17 (.BLUT(bypass_data_0_31__N_1012[16]), 
          .ALUT(bypass_data_0_31__N_882[16]), .C0(n37947), .Z(bypass_data_0[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i16 (.BLUT(bypass_data_0_31__N_1012[15]), 
          .ALUT(bypass_data_0_31__N_882[15]), .C0(n37947), .Z(bypass_data_0[15])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i8 (.BLUT(bypass_data_0_31__N_1012[7]), .ALUT(bypass_data_0_31__N_882[7]), 
          .C0(n37948), .Z(bypass_data_0[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i7 (.BLUT(bypass_data_0_31__N_1012[6]), .ALUT(bypass_data_0_31__N_882[6]), 
          .C0(n37952), .Z(bypass_data_0[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i6 (.BLUT(bypass_data_0_31__N_1012[5]), .ALUT(bypass_data_0_31__N_882[5]), 
          .C0(n36552), .Z(bypass_data_0[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i5 (.BLUT(bypass_data_0_31__N_1012[4]), .ALUT(bypass_data_0_31__N_882[4]), 
          .C0(n37950), .Z(bypass_data_0[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i4 (.BLUT(bypass_data_0_31__N_1012[3]), .ALUT(bypass_data_0_31__N_882[3]), 
          .C0(n37949), .Z(bypass_data_0[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i3 (.BLUT(bypass_data_0_31__N_1012[2]), .ALUT(bypass_data_0_31__N_882[2]), 
          .C0(n37953), .Z(bypass_data_0[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i2 (.BLUT(bypass_data_0_31__N_1012[1]), .ALUT(bypass_data_0_31__N_882[1]), 
          .C0(n37951), .Z(bypass_data_0[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i1 (.BLUT(n17974), .ALUT(bypass_data_1_31__N_914[0]), 
          .C0(n37940), .Z(bypass_data_1[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i1 (.BLUT(n17969), .ALUT(bypass_data_0_31__N_882[0]), 
          .C0(n37947), .Z(bypass_data_0[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_2_lut_rep_1095 (.A(branch_flushX_m), .B(dcache_refill_request), 
         .C(n41233), .D(cycles_5__N_2934), .Z(REF_CLK_c_enable_435)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1715[20] 1717[52])
    defparam i1_2_lut_rep_1095.init = 16'h0f0e;
    LUT4 operand_w_31__I_0_i3_3_lut (.A(operand_w[2]), .B(multiplier_result_w[2]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_690[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i3_3_lut.init = 16'hcaca;
    PFUMX bypass_data_1_31__I_0_i15 (.BLUT(bypass_data_1_31__N_1044[14]), 
          .ALUT(bypass_data_1_31__N_914[14]), .C0(n37944), .Z(bypass_data_1[14])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i14 (.BLUT(bypass_data_1_31__N_1044[13]), 
          .ALUT(bypass_data_1_31__N_914[13]), .C0(n37946), .Z(bypass_data_1[13])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i13 (.BLUT(bypass_data_1_31__N_1044[12]), 
          .ALUT(bypass_data_1_31__N_914[12]), .C0(n37942), .Z(bypass_data_1[12])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i12 (.BLUT(bypass_data_1_31__N_1044[11]), 
          .ALUT(bypass_data_1_31__N_914[11]), .C0(n37943), .Z(bypass_data_1[11])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i11 (.BLUT(bypass_data_1_31__N_1044[10]), 
          .ALUT(bypass_data_1_31__N_914[10]), .C0(n36614), .Z(bypass_data_1[10])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i10 (.BLUT(bypass_data_1_31__N_1044[9]), .ALUT(bypass_data_1_31__N_914[9]), 
          .C0(n37945), .Z(bypass_data_1[9])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i9 (.BLUT(bypass_data_1_31__N_1044[8]), .ALUT(bypass_data_1_31__N_914[8]), 
          .C0(n37941), .Z(bypass_data_1[8])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i15 (.BLUT(bypass_data_0_31__N_1012[14]), 
          .ALUT(bypass_data_0_31__N_882[14]), .C0(n37951), .Z(bypass_data_0[14])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i14 (.BLUT(bypass_data_0_31__N_1012[13]), 
          .ALUT(bypass_data_0_31__N_882[13]), .C0(n37953), .Z(bypass_data_0[13])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i13 (.BLUT(bypass_data_0_31__N_1012[12]), 
          .ALUT(bypass_data_0_31__N_882[12]), .C0(n37949), .Z(bypass_data_0[12])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i12 (.BLUT(bypass_data_0_31__N_1012[11]), 
          .ALUT(bypass_data_0_31__N_882[11]), .C0(n37950), .Z(bypass_data_0[11])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i11 (.BLUT(bypass_data_0_31__N_1012[10]), 
          .ALUT(bypass_data_0_31__N_882[10]), .C0(n36552), .Z(bypass_data_0[10])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i10 (.BLUT(bypass_data_0_31__N_1012[9]), 
          .ALUT(bypass_data_0_31__N_882[9]), .C0(n37952), .Z(bypass_data_0[9])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_13_i9 (.BLUT(bypass_data_0_31__N_1012[8]), .ALUT(bypass_data_0_31__N_882[8]), 
          .C0(n37948), .Z(bypass_data_0[8])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX i21 (.BLUT(logic_result_x[3]), .ALUT(n8), .C0(n37160), .Z(x_result[3]));
    PFUMX x_result_31__I_0_i32 (.BLUT(logic_result_x[31]), .ALUT(x_result_31__N_626[31]), 
          .C0(n36983), .Z(x_result[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 n10760_bdd_4_lut_33727 (.A(n41288), .B(n41391), .C(im[12]), .D(deba[12]), 
         .Z(n39327)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (D))) */ ;
    defparam n10760_bdd_4_lut_33727.init = 16'hec20;
    PFUMX x_result_31__I_0_i31 (.BLUT(logic_result_x[30]), .ALUT(x_result_31__N_626[30]), 
          .C0(n36971), .Z(x_result[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i30 (.BLUT(logic_result_x[29]), .ALUT(x_result_31__N_626[29]), 
          .C0(n36958), .Z(x_result[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i29 (.BLUT(logic_result_x[28]), .ALUT(x_result_31__N_626[28]), 
          .C0(n36945), .Z(x_result[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i28 (.BLUT(logic_result_x[27]), .ALUT(x_result_31__N_626[27]), 
          .C0(n36932), .Z(x_result[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX i34518 (.BLUT(logic_result_x[11]), .ALUT(n41750), .C0(n36724), 
          .Z(n41751));
    PFUMX x_result_31__I_0_i27 (.BLUT(logic_result_x[26]), .ALUT(x_result_31__N_626[26]), 
          .C0(n36919), .Z(x_result[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i26 (.BLUT(logic_result_x[25]), .ALUT(x_result_31__N_626[25]), 
          .C0(n36906), .Z(x_result[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i25 (.BLUT(logic_result_x[24]), .ALUT(x_result_31__N_626[24]), 
          .C0(n36893), .Z(x_result[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i24 (.BLUT(logic_result_x[23]), .ALUT(x_result_31__N_626[23]), 
          .C0(n36880), .Z(x_result[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i23 (.BLUT(logic_result_x[22]), .ALUT(x_result_31__N_626[22]), 
          .C0(n36867), .Z(x_result[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i22 (.BLUT(logic_result_x[21]), .ALUT(x_result_31__N_626[21]), 
          .C0(n36854), .Z(x_result[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i21 (.BLUT(logic_result_x[20]), .ALUT(x_result_31__N_626[20]), 
          .C0(n36841), .Z(x_result[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i20 (.BLUT(logic_result_x[19]), .ALUT(x_result_31__N_626[19]), 
          .C0(n36828), .Z(x_result[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i19 (.BLUT(logic_result_x[18]), .ALUT(x_result_31__N_626[18]), 
          .C0(n36815), .Z(x_result[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i18 (.BLUT(logic_result_x[17]), .ALUT(x_result_31__N_626[17]), 
          .C0(n36802), .Z(x_result[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i17 (.BLUT(logic_result_x[16]), .ALUT(x_result_31__N_626[16]), 
          .C0(n36789), .Z(x_result[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i16 (.BLUT(logic_result_x[15]), .ALUT(x_result_31__N_626[15]), 
          .C0(n36776), .Z(x_result[15])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i8 (.BLUT(logic_result_x[7]), .ALUT(x_result_31__N_626[7]), 
          .C0(n36686), .Z(x_result[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX i34435 (.BLUT(n41573), .ALUT(n41574), .C0(csr_x[3]), .Z(n41575));
    PFUMX x_result_31__I_0_i7 (.BLUT(logic_result_x[6]), .ALUT(x_result_31__N_626[6]), 
          .C0(n36673), .Z(x_result[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i6 (.BLUT(logic_result_x[5]), .ALUT(x_result_31__N_626[5]), 
          .C0(n36660), .Z(x_result[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i5 (.BLUT(logic_result_x[4]), .ALUT(x_result_31__N_626[4]), 
          .C0(n36647), .Z(x_result[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i3 (.BLUT(logic_result_x[2]), .ALUT(x_result_31__N_626[2]), 
          .C0(n36635), .Z(x_result[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i2 (.BLUT(logic_result_x[1]), .ALUT(x_result_31__N_626[1]), 
          .C0(n36623), .Z(x_result[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i1 (.BLUT(logic_result_x[0]), .ALUT(x_result_31__N_626[0]), 
          .C0(n36383), .Z(x_result[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX i34433 (.BLUT(n41570), .ALUT(n41571), .C0(csr_x[3]), .Z(n41572));
    PFUMX i34431 (.BLUT(n41567), .ALUT(n41568), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[6]));
    PFUMX i34429 (.BLUT(n41564), .ALUT(n41565), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[7]));
    PFUMX i34427 (.BLUT(n41561), .ALUT(n41562), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[8]));
    PFUMX i34515 (.BLUT(n41745), .ALUT(n41741), .C0(x_result_sel_csr_x), 
          .Z(n41746));
    PFUMX i34425 (.BLUT(n41558), .ALUT(n41559), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[9]));
    PFUMX i34423 (.BLUT(n41555), .ALUT(n41556), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[10]));
    PFUMX i34421 (.BLUT(n41552), .ALUT(n41553), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[11]));
    PFUMX i34513 (.BLUT(logic_result_x[10]), .ALUT(n41743), .C0(n36713), 
          .Z(n41744));
    PFUMX i34419 (.BLUT(n41549), .ALUT(n41550), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[12]));
    PFUMX i34417 (.BLUT(n41546), .ALUT(n41547), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[13]));
    PFUMX i34415 (.BLUT(n41543), .ALUT(n41544), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[14]));
    PFUMX i34413 (.BLUT(n41540), .ALUT(n41541), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[15]));
    PFUMX i34411 (.BLUT(n41537), .ALUT(n41538), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[16]));
    PFUMX i34409 (.BLUT(n41534), .ALUT(n41535), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[17]));
    PFUMX i34510 (.BLUT(n41738), .ALUT(n41734), .C0(x_result_sel_csr_x), 
          .Z(n41739));
    PFUMX i34407 (.BLUT(n41531), .ALUT(n41532), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[18]));
    PFUMX i34405 (.BLUT(n41528), .ALUT(n41529), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[19]));
    PFUMX i34403 (.BLUT(n41525), .ALUT(n41526), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[20]));
    LUT4 i1_4_lut_adj_642 (.A(n34556), .B(write_idx_w[4]), .C(n2_adj_6220), 
         .D(n41357), .Z(raw_w_1)) /* synthesis lut_function=(!((B (C+!(D))+!B (C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_642.init = 16'h0802;
    LUT4 i1_4_lut_adj_643 (.A(write_idx_w[3]), .B(n35591), .C(n41430), 
         .D(n41356), .Z(n34556)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_643.init = 16'h2010;
    PFUMX i34508 (.BLUT(logic_result_x[9]), .ALUT(n41736), .C0(n36702), 
          .Z(n41737));
    PFUMX i34401 (.BLUT(n41522), .ALUT(n41523), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[21]));
    PFUMX i34399 (.BLUT(n41519), .ALUT(n41520), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[22]));
    PFUMX i34397 (.BLUT(n41516), .ALUT(n41517), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[23]));
    PFUMX i34395 (.BLUT(n41513), .ALUT(n41514), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[24]));
    PFUMX i34503 (.BLUT(logic_result_x[8]), .ALUT(n41729), .C0(n36691), 
          .Z(n41730));
    PFUMX i34393 (.BLUT(n41510), .ALUT(n41511), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[25]));
    PFUMX i14156 (.BLUT(n19), .ALUT(n5780[7]), .C0(csr_x[2]), .Z(n3));
    PFUMX i34391 (.BLUT(n41507), .ALUT(n41508), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[26]));
    PFUMX i14160 (.BLUT(n18), .ALUT(n5780[6]), .C0(csr_x[2]), .Z(n5848[6]));
    PFUMX i34389 (.BLUT(n41504), .ALUT(n41505), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[27]));
    PFUMX i10 (.BLUT(n17), .ALUT(n5780[3]), .C0(csr_x[2]), .Z(n7));
    PFUMX i34387 (.BLUT(n41501), .ALUT(n41502), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[28]));
    PFUMX mux_2227_i32 (.BLUT(n5814[31]), .ALUT(n5780[31]), .C0(csr_x[2]), 
          .Z(n5848[31]));
    PFUMX mux_2227_i31 (.BLUT(n5814[30]), .ALUT(n5780[30]), .C0(csr_x[2]), 
          .Z(n5848[30]));
    PFUMX mux_2227_i30 (.BLUT(n5814[29]), .ALUT(n5780[29]), .C0(csr_x[2]), 
          .Z(n5848[29]));
    PFUMX mux_2227_i29 (.BLUT(n5814[28]), .ALUT(n5780[28]), .C0(csr_x[2]), 
          .Z(n5848[28]));
    LUT4 i30447_4_lut (.A(write_idx_w[2]), .B(n45103), .C(n41359), .D(n41355), 
         .Z(n35591)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i30447_4_lut.init = 16'h7bde;
    PFUMX i34385 (.BLUT(n41498), .ALUT(n41499), .C0(non_debug_exception_x), 
          .Z(branch_target_m_31__N_1167[29]));
    PFUMX mux_2227_i28 (.BLUT(n5814[27]), .ALUT(n5780[27]), .C0(csr_x[2]), 
          .Z(n5848[27]));
    PFUMX mux_2227_i27 (.BLUT(n5814[26]), .ALUT(n5780[26]), .C0(csr_x[2]), 
          .Z(n5848[26]));
    PFUMX mux_2227_i26 (.BLUT(n5814[25]), .ALUT(n5780[25]), .C0(csr_x[2]), 
          .Z(n5848[25]));
    PFUMX mux_2227_i25 (.BLUT(n5814[24]), .ALUT(n5780[24]), .C0(csr_x[2]), 
          .Z(n5848[24]));
    PFUMX mux_2227_i24 (.BLUT(n5814[23]), .ALUT(n5780[23]), .C0(csr_x[2]), 
          .Z(n5848[23]));
    PFUMX mux_2227_i23 (.BLUT(n5814[22]), .ALUT(n5780[22]), .C0(csr_x[2]), 
          .Z(n5848[22]));
    LUT4 i33156_rep_176_2_lut (.A(raw_x_1), .B(raw_m_1), .Z(n37940)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1529[10] 1534[36])
    defparam i33156_rep_176_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_644 (.A(n30245), .B(n35587), .C(n30012), .D(n5), 
         .Z(raw_m_1)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_644.init = 16'h0010;
    PFUMX mux_2227_i22 (.BLUT(n5814[21]), .ALUT(n5780[21]), .C0(csr_x[2]), 
          .Z(n5848[21]));
    PFUMX mux_2227_i21 (.BLUT(n5814[20]), .ALUT(n5780[20]), .C0(csr_x[2]), 
          .Z(n5848[20]));
    PFUMX mux_2227_i20 (.BLUT(n5814[19]), .ALUT(n5780[19]), .C0(csr_x[2]), 
          .Z(n5848[19]));
    LUT4 i33156_rep_180_2_lut (.A(raw_x_1), .B(raw_m_1), .Z(n37944)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1529[10] 1534[36])
    defparam i33156_rep_180_2_lut.init = 16'heeee;
    PFUMX mux_2227_i19 (.BLUT(n5814[18]), .ALUT(n5780[18]), .C0(csr_x[2]), 
          .Z(n5848[18]));
    PFUMX mux_2227_i18 (.BLUT(n5814[17]), .ALUT(n5780[17]), .C0(csr_x[2]), 
          .Z(n5848[17]));
    PFUMX mux_2227_i17 (.BLUT(n5814[16]), .ALUT(n5780[16]), .C0(csr_x[2]), 
          .Z(n5848[16]));
    PFUMX mux_2227_i16 (.BLUT(n5814[15]), .ALUT(n5780[15]), .C0(csr_x[2]), 
          .Z(n5848[15]));
    PFUMX mux_2227_i3 (.BLUT(n5814[2]), .ALUT(n5780[2]), .C0(csr_x[2]), 
          .Z(n5848[2]));
    LUT4 i33156_rep_182_2_lut (.A(raw_x_1), .B(raw_m_1), .Z(n37946)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1529[10] 1534[36])
    defparam i33156_rep_182_2_lut.init = 16'heeee;
    LUT4 i33156_rep_178_2_lut (.A(raw_x_1), .B(raw_m_1), .Z(n37942)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1529[10] 1534[36])
    defparam i33156_rep_178_2_lut.init = 16'heeee;
    PFUMX mux_2227_i2 (.BLUT(n5814[1]), .ALUT(n5780[1]), .C0(csr_x[2]), 
          .Z(n5848[1]));
    PFUMX w_result_31__I_0_i32 (.BLUT(w_result_31__N_690[31]), .ALUT(load_data_w[31]), 
          .C0(w_result_sel_load_w), .Z(w_result[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i33156_rep_179_2_lut (.A(raw_x_1), .B(raw_m_1), .Z(n37943)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1529[10] 1534[36])
    defparam i33156_rep_179_2_lut.init = 16'heeee;
    PFUMX w_result_31__I_0_i31 (.BLUT(w_result_31__N_690[30]), .ALUT(load_data_w[30]), 
          .C0(w_result_sel_load_w), .Z(w_result[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i30 (.BLUT(w_result_31__N_690[29]), .ALUT(load_data_w[29]), 
          .C0(w_result_sel_load_w), .Z(w_result[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i29 (.BLUT(w_result_31__N_690[28]), .ALUT(load_data_w[28]), 
          .C0(w_result_sel_load_w), .Z(w_result[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i28 (.BLUT(w_result_31__N_690[27]), .ALUT(load_data_w[27]), 
          .C0(w_result_sel_load_w), .Z(w_result[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i27 (.BLUT(w_result_31__N_690[26]), .ALUT(load_data_w[26]), 
          .C0(w_result_sel_load_w), .Z(w_result[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i26 (.BLUT(w_result_31__N_690[25]), .ALUT(load_data_w[25]), 
          .C0(w_result_sel_load_w), .Z(w_result[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i33156_2_lut (.A(raw_x_1), .B(raw_m_1), .Z(n36614)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1529[10] 1534[36])
    defparam i33156_2_lut.init = 16'heeee;
    PFUMX w_result_31__I_0_i25 (.BLUT(w_result_31__N_690[24]), .ALUT(load_data_w[24]), 
          .C0(w_result_sel_load_w), .Z(w_result[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i24 (.BLUT(w_result_31__N_690[23]), .ALUT(load_data_w[23]), 
          .C0(w_result_sel_load_w), .Z(w_result[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i33156_rep_181_2_lut (.A(raw_x_1), .B(raw_m_1), .Z(n37945)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1529[10] 1534[36])
    defparam i33156_rep_181_2_lut.init = 16'heeee;
    PFUMX w_result_31__I_0_i23 (.BLUT(w_result_31__N_690[22]), .ALUT(load_data_w[22]), 
          .C0(w_result_sel_load_w), .Z(w_result[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i22 (.BLUT(w_result_31__N_690[21]), .ALUT(load_data_w[21]), 
          .C0(w_result_sel_load_w), .Z(w_result[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i21 (.BLUT(w_result_31__N_690[20]), .ALUT(load_data_w[20]), 
          .C0(w_result_sel_load_w), .Z(w_result[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i20 (.BLUT(w_result_31__N_690[19]), .ALUT(load_data_w[19]), 
          .C0(w_result_sel_load_w), .Z(w_result[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i19 (.BLUT(w_result_31__N_690[18]), .ALUT(load_data_w[18]), 
          .C0(w_result_sel_load_w), .Z(w_result[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i18 (.BLUT(w_result_31__N_690[17]), .ALUT(load_data_w[17]), 
          .C0(w_result_sel_load_w), .Z(w_result[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i17 (.BLUT(w_result_31__N_690[16]), .ALUT(load_data_w[16]), 
          .C0(w_result_sel_load_w), .Z(w_result[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i33156_rep_177_2_lut (.A(raw_x_1), .B(raw_m_1), .Z(n37941)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1529[10] 1534[36])
    defparam i33156_rep_177_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_645 (.A(n35832), .B(n45099), .C(n33920), .D(n41354), 
         .Z(raw_w_0)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !((D)+!C)))) */ ;
    defparam i1_4_lut_adj_645.init = 16'h4010;
    PFUMX w_result_31__I_0_i8 (.BLUT(w_result_31__N_690[7]), .ALUT(load_data_w[7]), 
          .C0(w_result_sel_load_w), .Z(w_result[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i7 (.BLUT(w_result_31__N_690[6]), .ALUT(load_data_w[6]), 
          .C0(w_result_sel_load_w), .Z(w_result[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i6 (.BLUT(w_result_31__N_690[5]), .ALUT(load_data_w[5]), 
          .C0(w_result_sel_load_w), .Z(w_result[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i5 (.BLUT(w_result_31__N_690[4]), .ALUT(load_data_w[4]), 
          .C0(w_result_sel_load_w), .Z(w_result[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    lm32_shifter shifter (.\operand_1_x[4] (operand_1_x[4]), .\operand_1_x[3] (operand_1_x[3]), 
            .left_shift_result({left_shift_result[31], Open_9, Open_10, 
            Open_11, Open_12, Open_13, Open_14, Open_15, Open_16, 
            Open_17, Open_18, Open_19, Open_20, Open_21, Open_22, 
            Open_23, Open_24, Open_25, Open_26, Open_27, Open_28, 
            Open_29, Open_30, Open_31, Open_32, Open_33, Open_34, 
            Open_35, Open_36, Open_37, Open_38, Open_39}), .REF_CLK_c(REF_CLK_c), 
            .REF_CLK_c_enable_1624(REF_CLK_c_enable_1624), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .\operand_1_x[2] (operand_1_x[2]), .\operand_1_x[1] (\operand_1_x[1] ), 
            .\operand_1_x[0] (operand_1_x[0]), .operand_0_x({operand_0_x}), 
            .direction_x(direction_x), .direction_m(direction_m), .\condition_x[2] (condition_x[2]), 
            .REF_CLK_c_enable_1030(REF_CLK_c_enable_1030), .\left_shift_result[27] (left_shift_result[27]), 
            .\left_shift_result[25] (left_shift_result[25]), .\left_shift_result[21] (\left_shift_result[21] ), 
            .\left_shift_result[10] (\left_shift_result[10] ), .\left_shift_result[6] (left_shift_result[6]), 
            .\left_shift_result[4] (left_shift_result[4]), .\left_shift_result[0] (left_shift_result[0]), 
            .\shifter_result_m[1] (shifter_result_m[1]), .\shifter_result_m[2] (shifter_result_m[2]), 
            .\shifter_result_m[3] (shifter_result_m[3]), .\shifter_result_m[5] (shifter_result_m[5]), 
            .\shifter_result_m[7] (shifter_result_m[7]), .\shifter_result_m[8] (shifter_result_m[8]), 
            .\shifter_result_m[9] (shifter_result_m[9]), .\shifter_result_m[11] (shifter_result_m[11]), 
            .\shifter_result_m[12] (shifter_result_m[12]), .\shifter_result_m[13] (shifter_result_m[13]), 
            .\shifter_result_m[14] (shifter_result_m[14]), .\shifter_result_m[15] (shifter_result_m[15]), 
            .\shifter_result_m[16] (shifter_result_m[16]), .\shifter_result_m[17] (shifter_result_m[17]), 
            .\shifter_result_m[18] (shifter_result_m[18]), .\shifter_result_m[19] (shifter_result_m[19]), 
            .\shifter_result_m[20] (shifter_result_m[20]), .\shifter_result_m[22] (shifter_result_m[22]), 
            .\shifter_result_m[23] (shifter_result_m[23]), .\shifter_result_m[24] (shifter_result_m[24]), 
            .\shifter_result_m[26] (shifter_result_m[26]), .\shifter_result_m[28] (shifter_result_m[28]), 
            .\shifter_result_m[29] (shifter_result_m[29]), .\shifter_result_m[30] (shifter_result_m[30])) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1071[14] 1082[6])
    lm32_multiplier multiplier (.multiplier_result_w({multiplier_result_w}), 
            .REF_CLK_c(REF_CLK_c), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .GND_net(GND_net), .VCC_net(VCC_net), .operand_1_x({operand_1_x[31:2], 
            \operand_1_x[1] , operand_1_x[0]}), .operand_0_x({operand_0_x}), 
            .n45171(n45171)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1087[17] 1097[6])
    lm32_mc_arithmetic mc_arithmetic (.REF_CLK_c(REF_CLK_c), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .b({b}), .REF_CLK_c_enable_1366(REF_CLK_c_enable_1366), .d_result_1({d_result_1}), 
            .p({Open_40, \p[30] , \p[29] , \p[28] , \p[27] , \p[26] , 
            \p[25] , \p[24] , \p[23] , \p[22] , \p[21] , \p[20] , 
            \p[19] , \p[18] , \p[17] , \p[16] , \p[15] , \p[14] , 
            \p[13] , \p[12] , \p[11] , \p[10] , \p[9] , \p[8] , 
            \p[7] , \p[6] , \p[5] , \p[4] , \p[3] , \p[2] , \p[1] , 
            \p[0] }), .mc_result_x({mc_result_x}), .divide_by_zero_x(divide_by_zero_x), 
            .cycles_5__N_2934(cycles_5__N_2934), .\a[31] (\a[31] ), .GND_net(GND_net), 
            .VCC_net(VCC_net), .n32636(n32636), .n15(n15), .n41231(n41231), 
            .n45183(n45183), .t({t}), .d_result_0({d_result_0}), .n45181(n45181), 
            .n41216(n41216), .n41196(n41196), .q_d(q_d), .n32608(n32608), 
            .n41197(n41197), .n20863(n20863), .n32652(n32652)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1102[20] 1128[6])
    lm32_logic_op logic_op (.\condition_x[2] (condition_x[2]), .direction_x(direction_x), 
            .operand_0_x({operand_0_x}), .mc_result_x({mc_result_x}), .x_result_sel_mc_arith_x(x_result_sel_mc_arith_x), 
            .logic_result_x({logic_result_x}), .size_x({size_x}), .n36175(n36175), 
            .n36178(n36178), .n36184(n36184), .n36190(n36190), .n36193(n36193), 
            .n36196(n36196), .n36199(n36199), .n36223(n36223), .n36226(n36226), 
            .n36229(n36229), .n36232(n36232), .n36235(n36235), .n36238(n36238), 
            .n36241(n36241), .n36244(n36244), .n36247(n36247), .n36250(n36250), 
            .n36253(n36253), .n36256(n36256), .n36259(n36259), .n36262(n36262), 
            .n36265(n36265), .n36268(n36268), .n36283(n36283), .n36187(n36187)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1059[15] 1067[6])
    \lm32_load_store_unit(base_address=32'b0,limit=32'b01111111111111111)  load_store_unit (.n41402(n41402), 
            .\adder_result_x[1] (adder_result_x[1]), .\adder_result_x[0] (adder_result_x[0]), 
            .n45171(n45171), .n41283(n41283), .dcache_refill_request(dcache_refill_request), 
            .n41215(n41215), .REF_CLK_c(REF_CLK_c), .REF_CLK_c_enable_1235(REF_CLK_c_enable_1235), 
            .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), .size_x({size_x}), 
            .LM32D_DAT_O({LM32D_DAT_O}), .REF_CLK_c_enable_949(REF_CLK_c_enable_949), 
            .REF_CLK_c_enable_1221(REF_CLK_c_enable_1221), .SHAREDBUS_DAT_O({SHAREDBUS_DAT_O}), 
            .LM32D_SEL_O({LM32D_SEL_O}), .\LM32D_ADR_O[0] (\LM32D_ADR_O[0] ), 
            .size_w({Open_41, size_w[0]}), .\LM32D_CTI_O[0] (\LM32D_CTI_O[0] ), 
            .n38965(n38965), .\data_w[31] (data_w[31]), .\data_w[15] (data_w[15]), 
            .\operand_w[1] (operand_w[1]), .stall_wb_load(stall_wb_load), 
            .\data_w[30] (data_w[30]), .\data_w[29] (data_w[29]), .n30879(n30879), 
            .\data_w[28] (data_w[28]), .\data_w[27] (data_w[27]), .\data_w[26] (data_w[26]), 
            .\data_w[25] (data_w[25]), .\data_w[24] (data_w[24]), .store_operand_x({store_operand_x}), 
            .dcache_select_m(dcache_select_m), .dcache_select_x(dcache_select_x), 
            .wb_select_m(wb_select_m), .LM32D_STB_O(LM32D_STB_O), .n41388(n41388), 
            .\condition_x[2] (condition_x[2]), .LM32D_CYC_O(LM32D_CYC_O), 
            .REF_CLK_c_enable_1050(REF_CLK_c_enable_1050), .\load_data_w[16] (load_data_w[16]), 
            .\load_data_w[17] (load_data_w[17]), .\load_data_w[18] (load_data_w[18]), 
            .\load_data_w[19] (load_data_w[19]), .\load_data_w[20] (load_data_w[20]), 
            .\load_data_w[21] (load_data_w[21]), .\load_data_w[22] (load_data_w[22]), 
            .\load_data_w[23] (load_data_w[23]), .\load_data_w[24] (load_data_w[24]), 
            .\load_data_w[25] (load_data_w[25]), .\load_data_w[26] (load_data_w[26]), 
            .\load_data_w[27] (load_data_w[27]), .\load_data_w[28] (load_data_w[28]), 
            .\load_data_w[29] (load_data_w[29]), .\load_data_w[30] (load_data_w[30]), 
            .\load_data_w[31] (load_data_w[31]), .LM32D_WE_O(LM32D_WE_O), 
            .REF_CLK_c_enable_1234(REF_CLK_c_enable_1234), .n12404(n12404), 
            .wb_load_complete(wb_load_complete), .REF_CLK_c_enable_1236(REF_CLK_c_enable_1236), 
            .n12400(n12400), .n21(n21), .\LM32D_ADR_O[1] (\LM32D_ADR_O[1] ), 
            .\LM32D_ADR_O[2] (\LM32D_ADR_O[2] ), .\next_cycle_type[2] (\next_cycle_type[2] ), 
            .\LM32D_ADR_O[4] (\LM32D_ADR_O[4] ), .\LM32D_ADR_O[5] (\LM32D_ADR_O[5] ), 
            .\d_adr_o_31__N_2278[5] (\d_adr_o_31__N_2278[5] ), .\LM32D_ADR_O[6] (\LM32D_ADR_O[6] ), 
            .\LM32D_ADR_O[7] (\LM32D_ADR_O[7] ), .\LM32D_ADR_O[8] (\LM32D_ADR_O[8] ), 
            .\LM32D_ADR_O[9] (\LM32D_ADR_O[9] ), .\d_adr_o_31__N_2278[9] (\d_adr_o_31__N_2278[9] ), 
            .\LM32D_ADR_O[10] (\LM32D_ADR_O[10] ), .\d_adr_o_31__N_2278[10] (\d_adr_o_31__N_2278[10] ), 
            .\LM32D_ADR_O[11] (\LM32D_ADR_O[11] ), .\LM32D_ADR_O[12] (\LM32D_ADR_O[12] ), 
            .\LM32D_ADR_O[13] (\LM32D_ADR_O[13] ), .\LM32D_ADR_O[14] (\LM32D_ADR_O[14] ), 
            .\LM32D_ADR_O[15] (\LM32D_ADR_O[15] ), .\LM32D_ADR_O[16] (\LM32D_ADR_O[16] ), 
            .\LM32D_ADR_O[17] (\LM32D_ADR_O[17] ), .\LM32D_ADR_O[18] (\LM32D_ADR_O[18] ), 
            .\LM32D_ADR_O[19] (\LM32D_ADR_O[19] ), .\LM32D_ADR_O[20] (\LM32D_ADR_O[20] ), 
            .\LM32D_ADR_O[21] (\LM32D_ADR_O[21] ), .\LM32D_ADR_O[22] (\LM32D_ADR_O[22] ), 
            .\LM32D_ADR_O[23] (\LM32D_ADR_O[23] ), .\LM32D_ADR_O[24] (\LM32D_ADR_O[24] ), 
            .\LM32D_ADR_O[25] (\LM32D_ADR_O[25] ), .\d_adr_o_31__N_2278[25] (d_adr_o_31__N_2278[25]), 
            .\LM32D_ADR_O[26] (\LM32D_ADR_O[26] ), .\LM32D_ADR_O[27] (\LM32D_ADR_O[27] ), 
            .\d_adr_o_31__N_2278[27] (d_adr_o_31__N_2278[27]), .\LM32D_ADR_O[28] (\LM32D_ADR_O[28] ), 
            .\LM32D_ADR_O[29] (\LM32D_ADR_O[29] ), .\LM32D_ADR_O[30] (\LM32D_ADR_O[30] ), 
            .\LM32D_ADR_O[31] (\LM32D_ADR_O[31] ), .REF_CLK_c_enable_1299(REF_CLK_c_enable_1299), 
            .REF_CLK_c_enable_1304(REF_CLK_c_enable_1304), .\data_w[8] (data_w[8]), 
            .\data_w[9] (data_w[9]), .\data_w[10] (data_w[10]), .\data_w[11] (data_w[11]), 
            .\data_w[12] (data_w[12]), .\data_w[13] (data_w[13]), .\data_w[14] (data_w[14]), 
            .\operand_w[0] (operand_w[0]), .dcache_refilling(dcache_refilling), 
            .n41387(n41387), .n20639(n20639), .n41380(n41380), .locked_N_493(locked_N_493), 
            .operand_m({operand_m[31:11], \operand_m[10] , \operand_m[9] , 
            operand_m[8:6], \operand_m[5] , operand_m[4:0]}), .n41217(n41217), 
            .exception_m(exception_m), .n41232(n41232), .n30070(n30070), 
            .n35745(n35745), .n41233(n41233), .n9(n9), .\load_data_w[6] (load_data_w[6]), 
            .n41144(n41144), .n41145(n41145), .n41156(n41156), .n41157(n41157), 
            .n41140(n41140), .n41141(n41141), .n41164(n41164), .n41165(n41165), 
            .n41160(n41160), .n41161(n41161), .\load_data_w[7] (load_data_w[7]), 
            .\load_data_w[5] (load_data_w[5]), .\load_data_w[4] (load_data_w[4]), 
            .n41148(n41148), .n41149(n41149), .\load_data_w[3] (load_data_w[3]), 
            .n41152(n41152), .n41153(n41153), .\load_data_w[2] (load_data_w[2]), 
            .n41136(n41136), .n41137(n41137), .\load_data_w[1] (load_data_w[1]), 
            .\load_data_w[0] (load_data_w[0]), .icache_refill_request(icache_refill_request), 
            .n41435(n41435), .branch_taken_m(branch_taken_m), .n41203(n41203), 
            .valid_d(valid_d), .q_d(q_d), .n32652(n32652), .\d_adr_o_31__N_2278[3] (d_adr_o_31__N_2278[3]), 
            .\d_adr_o_31__N_2278[2] (d_adr_o_31__N_2278[2]), .dcache_restart_request(dcache_restart_request), 
            .n45183(n45183), .state({\state[2] , state_adj_6256[1], \state[0] }), 
            .flush_set({flush_set}), .flush_set_8__N_2513({flush_set_8__N_2513}), 
            .\dcache_refill_address[5] (\dcache_refill_address[5] ), .\dcache_refill_address[9] (\dcache_refill_address[9] ), 
            .\dcache_refill_address[10] (\dcache_refill_address[10] ), .\dcache_refill_address[25] (dcache_refill_address[25]), 
            .\dcache_refill_address[27] (dcache_refill_address[27]), .n41284(n41284), 
            .icache_restart_request(icache_restart_request), .n19852(n19852), 
            .valid_a(valid_a), .n30107(n30107), .n9304(n9304), .\state[2]_adj_192 (state[2]), 
            .n41187(n41187), .n41196(n41196), .n31996(n31996), .n45175(n45175), 
            .way_match_0__N_2007(way_match_0__N_2007), .valid_f(valid_f), 
            .dflush_m(dflush_m), .n41178(n41178), .n36389(n36389), .n37914(n37914), 
            .n37915(n37915), .n37919(n37919), .n37917(n37917), .n37916(n37916), 
            .n37918(n37918), .n41(n41), .restart_request_N_1998(restart_request_N_1998), 
            .n15(n15), .n41172(n41172), .n32278(n32278), .\tmem_write_address[1] (\tmem_write_address[1] ), 
            .\tmem_write_address[5] (\tmem_write_address[5] ), .\tmem_write_address[6] (\tmem_write_address[6] ), 
            .n7502({n7502}), .VCC_net(VCC_net), .GND_net(GND_net), .\genblk1.ra ({\genblk1.ra_adj_6257 }), 
            .\dmem_write_address[3] (\dmem_write_address[3] ), .\dmem_write_address[7] (\dmem_write_address[7] ), 
            .\dmem_write_address[8] (\dmem_write_address[8] ), .n7388({n7388}), 
            .n7322({n7322}), .n7256({n7256}), .n7204(n7204), .n7190({n7190}), 
            .n7206(n7206), .n7208(n7208), .\genblk1.ra_adj_202 ({\genblk1.ra }), 
            .n7224(n7224), .n7222(n7222), .n7220(n7220), .n7356(n7356), 
            .n7354(n7354), .n7352(n7352), .n7350(n7350), .n7348(n7348), 
            .n7346(n7346), .n7344(n7344), .n7342(n7342), .n7340(n7340), 
            .n7338(n7338), .n7336(n7336), .n7218(n7218), .n7290(n7290), 
            .n7288(n7288), .n7286(n7286), .n7284(n7284), .n7216(n7216), 
            .n7282(n7282), .n7280(n7280), .n7278(n7278), .n7214(n7214), 
            .n7276(n7276), .n7274(n7274), .n7272(n7272), .n7212(n7212), 
            .n7270(n7270), .n7210(n7210)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(984[5] 1043[6])
    lm32_jtag jtag (.jtag_reg_q({jtag_reg_q}), .jtag_reg_d_7__N_515(jtag_reg_d_7__N_515), 
            .jtag_reg_d({jtag_reg_d}), .REF_CLK_c(REF_CLK_c), .REF_CLK_c_enable_1373(REF_CLK_c_enable_1373), 
            .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), .n4626({n4626}), 
            .rx_toggle_r_r(rx_toggle_r_r), .rx_toggle_r_r_r(rx_toggle_r_r_r), 
            .uart_tx_byte({uart_tx_byte}), .\operand_1_x[0] (operand_1_x[0]), 
            .\jrx_csr_read_data[0] (jrx_csr_read_data[0]), .jrx_csr_read_data_8__N_3304(jrx_csr_read_data_8__N_3304), 
            .jtag_break(jtag_break), .reset_exception(reset_exception), 
            .\jtag_reg_addr_d[0] (\jtag_reg_addr_d[0] ), .\jtag_reg_addr_d[1] (\jtag_reg_addr_d[1] ), 
            .jtag_update_N_3371(jtag_update_N_3371), .\operand_1_x[1] (\operand_1_x[1] ), 
            .\operand_1_x[2] (operand_1_x[2]), .\operand_1_x[3] (operand_1_x[3]), 
            .\operand_1_x[4] (operand_1_x[4]), .\operand_1_x[5] (operand_1_x[5]), 
            .\operand_1_x[6] (operand_1_x[6]), .\operand_1_x[7] (operand_1_x[7]), 
            .\jrx_csr_read_data[1] (jrx_csr_read_data[1]), .\jrx_csr_read_data[2] (jrx_csr_read_data[2]), 
            .\jrx_csr_read_data[3] (jrx_csr_read_data[3]), .\jrx_csr_read_data[4] (jrx_csr_read_data[4]), 
            .\jrx_csr_read_data[5] (jrx_csr_read_data[5]), .\jrx_csr_read_data[6] (jrx_csr_read_data[6]), 
            .\jrx_csr_read_data[7] (jrx_csr_read_data[7]), .n41232(n41232), 
            .n4(n4), .n41233(n41233), .n34542(n34542), .\jtag_reg_addr_q[1] (\jtag_reg_addr_q[1] ), 
            .n30162(n30162), .n43(n43), .n33932(n33932), .n29834(n29834), 
            .n34464(n34464)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1163[11] 1208[6])
    lm32_interrupt interrupt (.csr_x({csr_x}), .n41288(n41288), .im({Open_42, 
            Open_43, Open_44, Open_45, Open_46, Open_47, Open_48, 
            Open_49, Open_50, Open_51, Open_52, Open_53, Open_54, 
            Open_55, Open_56, Open_57, Open_58, Open_59, Open_60, 
            Open_61, Open_62, Open_63, Open_64, Open_65, Open_66, 
            Open_67, Open_68, Open_69, Open_70, Open_71, Open_72, 
            im[0]}), .REF_CLK_c(REF_CLK_c), .REF_CLK_c_enable_1335(REF_CLK_c_enable_1335), 
            .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), .operand_1_x({operand_1_x[31:2], 
            \operand_1_x[1] , operand_1_x[0]}), .n41308(n41308), .n4354(n4323[1]), 
            .bie(bie), .REF_CLK_c_enable_391(REF_CLK_c_enable_391), .n36337(n36337), 
            .n9401(n9401), .ie(ie), .\im[2] (im[2]), .\im[3] (im[3]), 
            .\im[4] (im[4]), .\im[5] (im[5]), .\im[6] (im[6]), .\im[7] (im[7]), 
            .\im[8] (im[8]), .\im[9] (im[9]), .\im[10] (im[10]), .\im[11] (im[11]), 
            .\im[12] (im[12]), .\im[13] (im[13]), .\im[14] (im[14]), .\im[15] (im[15]), 
            .\im[16] (im[16]), .\im[17] (im[17]), .\im[18] (im[18]), .\im[19] (im[19]), 
            .\im[20] (im[20]), .\im[21] (im[21]), .\im[22] (im[22]), .\im[23] (im[23]), 
            .\im[24] (im[24]), .\im[25] (im[25]), .\im[26] (im[26]), .\im[27] (im[27]), 
            .\im[28] (im[28]), .\im[29] (im[29]), .\im[30] (im[30]), .\im[31] (im[31]), 
            .\ip[1] (ip[1]), .n32134(n32134), .store_x(store_x), .n32132(n32132), 
            .n41313(n41313), .n41393(n41393), .n41391(n41391), .n31825(n31825), 
            .n11934(n11934), .n45175(n45175), .branch_flushX_m(branch_flushX_m), 
            .n35639(n35639), .dcache_refill_request(dcache_refill_request), 
            .n35022(n35022), .eret_q_x(eret_q_x), .n34986(n34986), .n35030(n35030), 
            .valid_w(valid_w), .non_debug_exception_w(non_debug_exception_w), 
            .debug_exception_w(debug_exception_w), .n41240(n41240), .n41394(n41394), 
            .eret_x(eret_x), .bret_x(bret_x), .n41400(n41400), .n34542(n34542), 
            .valid_x(valid_x), .n20581(n20581), .n41232(n41232), .n34942(n34942), 
            .SPI_INT_O_N_4422(SPI_INT_O_N_4422), .SPI_INT_O_N_4417(SPI_INT_O_N_4417), 
            .SPI_INT_O_N_4421(SPI_INT_O_N_4421), .n31334(n31334), .n41183(n41183), 
            .n41401(n41401), .n41317(n41317), .n41413(n41413), .n34898(n34898), 
            .n41416(n41416), .LM32D_CYC_O(LM32D_CYC_O), .n33946(n33946)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1133[16] 1158[6])
    \lm32_instruction_unit(base_address=32'b0,limit=32'b01111111111111111)  instruction_unit (.\genblk1.wait_one_tick_done (\genblk1.wait_one_tick_done ), 
            .n6781(n6781), .n41208(n41208), .n6764(n6764), .n6769(n6769), 
            .n6749(n6749), .REF_CLK_c(REF_CLK_c), .stall_a(stall_a), .way_match_0__N_2007(way_match_0__N_2007), 
            .bus_error_f_N_1884(bus_error_f_N_1884), .n41410(n41410), .n13990(n13990), 
            .n32216(n32216), .n45075(n45075), .n41244(n41244), .n41419(n41419), 
            .n41295(n41295), .n41248(n41248), .n30216(n30216), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .VCC_net(VCC_net), .n41178(n41178), .\LM32I_CTI_O[0] (\LM32I_CTI_O[0] ), 
            .REF_CLK_c_enable_97(REF_CLK_c_enable_97), .n30900(n30900), 
            .pc_d({pc_d}), .REF_CLK_c_enable_1178(REF_CLK_c_enable_1178), 
            .pc_f({pc_f}), .pc_x({pc_x}), .REF_CLK_c_enable_1624(REF_CLK_c_enable_1624), 
            .pc_m({pc_m}), .REF_CLK_c_enable_1235(REF_CLK_c_enable_1235), 
            .REF_CLK_c_enable_1131(REF_CLK_c_enable_1131), .SHAREDBUS_DAT_O({SHAREDBUS_DAT_O}), 
            .n6760(n6760), .n6765(n6765), .n31717(n31717), .n45105(n45105), 
            .n6771(n6771), .n73(n73), .n41461(n41461), .n41228(n41228), 
            .n41365(n41365), .n41361(n41361), .scall_d(scall_d), .n41437(n41437), 
            .n6778(n6778), .n6780(n6780), .n31542(n31542), .n6768(n6768), 
            .n32910(n32910), .n6779(n6779), .n10(n10), .n6777(n6777), 
            .n6775(n6775), .branch_taken_m(branch_taken_m), .icache_refill_request(icache_refill_request), 
            .\next_cycle_type[2] (\next_cycle_type[2]_adj_203 ), .n45080(n45080), 
            .n41390(n41390), .n5223(n5223), .n37955(n37955), .n37956(n37956), 
            .n37954(n37954), .n41345(n41345), .n41250(n41250), .n41251(n41251), 
            .n41279(n41279), .\LM32I_ADR_O[2] (\LM32I_ADR_O[2] ), .n45079(n45079), 
            .\reg_12[2] (\reg_12[2] ), .n2(n2), .\reg_12[12] (\reg_12[12] ), 
            .n40677(n40677), .\reg_12[29] (\reg_12[29] ), .n2_adj_149(n2_adj_204), 
            .\reg_12[3] (\reg_12[3] ), .n2_adj_150(n2_adj_205), .\reg_12[6] (\reg_12[6] ), 
            .n2_adj_151(n2_adj_206), .\reg_12[4] (\reg_12[4] ), .n2_adj_152(n2_adj_207), 
            .\reg_12[14] (\reg_12[14] ), .n2_adj_153(n2_adj_208), .n30241(n30241), 
            .n31750(n31750), .n31955(n31955), .n41429(n41429), .\reg_12[22] (\reg_12[22] ), 
            .n2_adj_154(n2_adj_209), .\reg_12[13] (\reg_12[13] ), .n2_adj_155(n2_adj_210), 
            .\reg_12[21] (\reg_12[21] ), .n2_adj_156(n2_adj_211), .\reg_12[28] (\reg_12[28] ), 
            .n2_adj_157(n2_adj_212), .\reg_12[11] (\reg_12[11] ), .n2_adj_158(n2_adj_213), 
            .\reg_12[18] (\reg_12[18] ), .n2_adj_159(n2_adj_214), .\reg_12[25] (\reg_12[25] ), 
            .n2_adj_160(n2_adj_215), .\reg_12[9] (\reg_12[9] ), .n2_adj_161(n2_adj_216), 
            .\reg_12[17] (\reg_12[17] ), .n2_adj_162(n2_adj_217), .\reg_12[24] (\reg_12[24] ), 
            .n2_adj_163(n2_adj_218), .\reg_12[7] (\reg_12[7] ), .n2_adj_164(n2_adj_219), 
            .\reg_12[15] (\reg_12[15] ), .n2_adj_165(n2_adj_220), .n41382(n41382), 
            .n45183(n45183), .n6770(n6770), .n6589(n6589), .n6584(n6584), 
            .n37179(n37179), .\write_idx_x[0] (write_idx_x[0]), .n35751(n35751), 
            .n35860(n35860), .n6439(n6439), .n6434(n6434), .n37177(n37177), 
            .n6599(n6599), .n6594(n6594), .n37180(n37180), .n6629(n6629), 
            .n6624(n6624), .n37183(n37183), .n6579(n6579), .n6574(n6574), 
            .n37178(n37178), .n6429(n6429), .n6424(n6424), .n37176(n37176), 
            .n45103(n45103), .n35687(n35687), .n35832(n35832), .n6609(n6609), 
            .n6604(n6604), .n37181(n37181), .n6619(n6619), .n6614(n6614), 
            .n37182(n37182), .n37185(n37185), .n37184(n37184), .n37188(n37188), 
            .n37187(n37187), .n37186(n37186), .n37189(n37189), .n7603(n7603), 
            .n7571(n7571), .n7609({n7609}), .n7607(n7607), .n7575(n7575), 
            .n7606(n7606), .n7574(n7574), .bus_error_d(bus_error_d), .n7604(n7604), 
            .n7572(n7572), .n7605(n7605), .n7573(n7573), .n7608(n7608), 
            .n7576(n7576), .n7602(n7602), .n7570(n7570), .\selected_1__N_354[0] (\selected_1__N_354[0] ), 
            .n7601(n7601), .n7569(n7569), .n7600(n7600), .n7568(n7568), 
            .n7599(n7599), .n7567(n7567), .n7598(n7598), .n7566(n7566), 
            .n7597(n7597), .n7565(n7565), .n7596(n7596), .n7564(n7564), 
            .n7595(n7595), .n7563(n7563), .n7594(n7594), .n7562(n7562), 
            .n7593(n7593), .n7561(n7561), .n7592(n7592), .n7560(n7560), 
            .n7584(n7584), .n7552(n7552), .n7583(n7583), .n7551(n7551), 
            .n7582(n7582), .n7550(n7550), .n7581(n7581), .n7549(n7549), 
            .n7580(n7580), .n7548(n7548), .n7579(n7579), .n7547(n7547), 
            .n7578(n7578), .n7546(n7546), .n7577(n7577), .n7545(n7545), 
            .n6750(n6750), .n7591(n7591), .n7559(n7559), .n7590(n7590), 
            .n7558(n7558), .n7589(n7589), .n7557(n7557), .n7588(n7588), 
            .n7556(n7556), .n7587(n7587), .n7555(n7555), .n7586(n7586), 
            .n7554(n7554), .n7585(n7585), .n7553(n7553), .n4(n4_adj_6193), 
            .\write_idx_x[3] (write_idx_x[3]), .n32116(n32116), .n41430(n41430), 
            .\write_idx_w[3] (write_idx_w[3]), .n33920(n33920), .n37501(n37501), 
            .n37500(n37500), .n37502(n37502), .n37499(n37499), .n37498(n37498), 
            .n37497(n37497), .n37496(n37496), .n6751(n6751), .n6752(n6752), 
            .n6753(n6753), .n6754(n6754), .n6755(n6755), .n6756(n6756), 
            .n6757(n6757), .n6758(n6758), .n6759(n6759), .n6761(n6761), 
            .n6762(n6762), .n6763(n6763), .n6766(n6766), .n6767(n6767), 
            .n6776(n6776), .n40094(n40094), .n37495(n37495), .n7672(n7672), 
            .n7640(n7640), .n7677({n7677}), .n7673(n7673), .n7641(n7641), 
            .\write_idx_x[4] (write_idx_x[4]), .n32260(n32260), .n32262(n32262), 
            .n41312(n41312), .n41296(n41296), .n34(n34), .n7674(n7674), 
            .n7642(n7642), .n7675(n7675), .n7643(n7643), .n7676(n7676), 
            .n7644(n7644), .n7671(n7671), .n7639(n7639), .n7670(n7670), 
            .n7638(n7638), .n7669(n7669), .n7637(n7637), .n7668(n7668), 
            .n7636(n7636), .n7667(n7667), .n7635(n7635), .n7666(n7666), 
            .n7634(n7634), .n7665(n7665), .n7633(n7633), .n7664(n7664), 
            .n7632(n7632), .n7663(n7663), .n7631(n7631), .n7662(n7662), 
            .n7630(n7630), .n7661(n7661), .n7629(n7629), .n7660(n7660), 
            .n7628(n7628), .n36(n36), .n7652(n7652), .n7620(n7620), 
            .n7651(n7651), .n7619(n7619), .n7650(n7650), .n7618(n7618), 
            .n7649(n7649), .n7617(n7617), .n37(n37), .n7648(n7648), 
            .n7616(n7616), .n7647(n7647), .n7615(n7615), .n7646(n7646), 
            .n7614(n7614), .n7645(n7645), .n7613(n7613), .n7659(n7659), 
            .n7627(n7627), .n7658(n7658), .n7626(n7626), .n7657(n7657), 
            .n7625(n7625), .n7656(n7656), .n7624(n7624), .n7655(n7655), 
            .n7623(n7623), .n7654(n7654), .n7622(n7622), .n7653(n7653), 
            .n7621(n7621), .n30012(n30012), .\write_idx_m[2] (write_idx_m[2]), 
            .n31976(n31976), .n37504(n37504), .n37503(n37503), .n37507(n37507), 
            .n37506(n37506), .n37505(n37505), .n37508(n37508), .n41364(n41364), 
            .n41363(n41363), .n30820(n30820), .n11834(n11834), .n41216(n41216), 
            .n32356(n32356), .n41281(n41281), .n41367(n41367), .n41441(n41441), 
            .n41229(n41229), .n41227(n41227), .n41319(n41319), .w_result_sel_mul_d(w_result_sel_mul_d), 
            .n41381(n41381), .n41451(n41451), .REF_CLK_c_enable_1030(REF_CLK_c_enable_1030), 
            .n45106(n45106), .REF_CLK_c_enable_1042(REF_CLK_c_enable_1042), 
            .REF_CLK_c_enable_1050(REF_CLK_c_enable_1050), .REF_CLK_c_enable_1299(REF_CLK_c_enable_1299), 
            .\LM32I_ADR_O[4] (\LM32I_ADR_O[4] ), .\LM32I_ADR_O[5] (\LM32I_ADR_O[5] ), 
            .\LM32I_ADR_O[6] (\LM32I_ADR_O[6] ), .\LM32I_ADR_O[7] (\LM32I_ADR_O[7] ), 
            .\LM32I_ADR_O[8] (\LM32I_ADR_O[8] ), .\LM32I_ADR_O[9] (\LM32I_ADR_O[9] ), 
            .\LM32I_ADR_O[10] (\LM32I_ADR_O[10] ), .\LM32I_ADR_O[11] (\LM32I_ADR_O[11] ), 
            .\LM32I_ADR_O[12] (\LM32I_ADR_O[12] ), .\LM32I_ADR_O[13] (\LM32I_ADR_O[13] ), 
            .\LM32I_ADR_O[14] (\LM32I_ADR_O[14] ), .\LM32I_ADR_O[15] (\LM32I_ADR_O[15] ), 
            .\LM32I_ADR_O[16] (\LM32I_ADR_O[16] ), .\LM32I_ADR_O[17] (\LM32I_ADR_O[17] ), 
            .\LM32I_ADR_O[18] (\LM32I_ADR_O[18] ), .\LM32I_ADR_O[19] (\LM32I_ADR_O[19] ), 
            .\LM32I_ADR_O[20] (\LM32I_ADR_O[20] ), .\LM32I_ADR_O[21] (\LM32I_ADR_O[21] ), 
            .\LM32I_ADR_O[22] (\LM32I_ADR_O[22] ), .\LM32I_ADR_O[23] (\LM32I_ADR_O[23] ), 
            .\LM32I_ADR_O[24] (\LM32I_ADR_O[24] ), .\LM32I_ADR_O[25] (\LM32I_ADR_O[25] ), 
            .\LM32I_ADR_O[26] (\LM32I_ADR_O[26] ), .\LM32I_ADR_O[27] (\LM32I_ADR_O[27] ), 
            .\LM32I_ADR_O[28] (\LM32I_ADR_O[28] ), .\LM32I_ADR_O[29] (\LM32I_ADR_O[29] ), 
            .\LM32I_ADR_O[30] (\LM32I_ADR_O[30] ), .\LM32I_ADR_O[31] (\LM32I_ADR_O[31] ), 
            .REF_CLK_c_enable_1425(REF_CLK_c_enable_1425), .n41285(n41285), 
            .n30888(n30888), .n41350(n41350), .n41351(n41351), .n41247(n41247), 
            .n41348(n41348), .\instruction_d[11] (instruction_d[11]), .\instruction_d[12] (instruction_d[12]), 
            .\instruction_d[13] (instruction_d[13]), .\instruction_d[14] (instruction_d[14]), 
            .n41352(n41352), .n41353(n41353), .n41354(n41354), .\write_idx_m[1] (write_idx_m[1]), 
            .n2_adj_166(n2_c), .\write_idx_x[1] (write_idx_x[1]), .n2_adj_167(n2_adj_6194), 
            .n41355(n41355), .n41356(n41356), .n41357(n41357), .\write_idx_m[4] (write_idx_m[4]), 
            .n5(n5), .n41358(n41358), .n45099(n45099), .n2_adj_168(n2_adj_6220), 
            .n41282(n41282), .n41359(n41359), .n10475(n10475), .n41366(n41366), 
            .n41368(n41368), .n41369(n41369), .n41370(n41370), .n41371(n41371), 
            .n41372(n41372), .pc_a_31__N_1720({pc_a_31__N_1720}), .n41373(n41373), 
            .n41374(n41374), .n41375(n41375), .n41376(n41376), .n41377(n41377), 
            .n41179(n41179), .\extended_immediate[31] (extended_immediate[31]), 
            .n2_adj_169(n2_adj_6241), .n41291(n41291), .n2_adj_170(n2_adj_6219), 
            .n2_adj_171(n2_adj_6242), .n2_adj_172(n2_adj_6218), .n2_adj_173(n2_adj_6243), 
            .n2_adj_174(n2_adj_6217), .n2_adj_175(n2_adj_6244), .n2_adj_176(n2_adj_6216), 
            .n6028(n6028), .n41232(n41232), .n35032(n35032), .n12412(n12412), 
            .dcache_refilling(dcache_refilling), .dcache_refill_request(dcache_refill_request), 
            .dcache_restart_request(dcache_restart_request), .n949({n949}), 
            .n32220(n32220), .locked_N_493(locked_N_493), .n40093(n40093), 
            .write_idx_d({write_idx_d}), .n41380(n41380), .LM32D_CYC_O(LM32D_CYC_O), 
            .n30879(n30879), .n10485(n10485), .n31519(n31519), .selected({selected}), 
            .m_result_sel_shift_d(m_result_sel_shift_d), .n30058(n30058), 
            .n41362(n41362), .LM32D_WE_O(LM32D_WE_O), .\LM32D_ADR_O[1] (\LM32D_ADR_O[1] ), 
            .n41452(n41452), .n41241(n41241), .n37918(n37918), .n37916(n37916), 
            .n37917(n37917), .n37919(n37919), .n37915(n37915), .n37914(n37914), 
            .n36389(n36389), .flush_set({flush_set_adj_231}), .icache_restart_request(icache_restart_request), 
            .restart_request_N_1998(restart_request_N_1998), .icache_refilling(icache_refilling), 
            .\state[2] (state[2]), .n41196(n41196), .n15(n15), .q_d(q_d), 
            .n45175(n45175), .valid_x_N_1285(valid_x_N_1285), .n32278(n32278), 
            .n10_adj_177(n10_adj_6254), .n32264(n32264), .n41203(n41203), 
            .n41408(n41408), .flush_set_8__N_1953({flush_set_8__N_1953}), 
            .n9304(n9304), .n41(n41), .n41187(n41187), .branch_target_d({branch_target_d}), 
            .n157({n157}), .n31996(n31996), .cycles_5__N_2934(cycles_5__N_2934), 
            .REF_CLK_c_enable_1366(REF_CLK_c_enable_1366), .REF_CLK_c_enable_1622(REF_CLK_c_enable_1622), 
            .n41172(n41172), .n32618(n32618), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(804[5] 896[6])
    \lm32_debug(watchpoints=32'b0)  hw_debug (.dc_re(dc_re), .REF_CLK_c(REF_CLK_c), 
            .REF_CLK_c_enable_388(REF_CLK_c_enable_388), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .n36336(n36336)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1216[5] 1249[6])
    lm32_decoder decoder (.n45106(n45106), .n41365(n41365), .n41362(n41362), 
            .n11807(n11807), .n41244(n41244), .n41247(n41247), .n6028(n6028), 
            .n41295(n41295), .n45075(n45075), .VCC_net(VCC_net), .n6777(n6777), 
            .n11834(n11834), .n41228(n41228), .n20863(n20863), .n41198(n41198), 
            .n30058(n30058), .n41381(n41381), .\bypass_data_0[0] (bypass_data_0[0]), 
            .\d_result_0[0] (d_result_0[0]), .\bypass_data_0[1] (bypass_data_0[1]), 
            .\d_result_0[1] (d_result_0[1]), .n41363(n41363), .n31717(n31717), 
            .bret_d(bret_d), .n6779(n6779), .\genblk1.wait_one_tick_done (\genblk1.wait_one_tick_done ), 
            .n6780(n6780), .n6770(n6770), .n6781(n6781), .n6775(n6775), 
            .n6776(n6776), .n10475(n10475), .n41382(n41382), .n6778(n6778), 
            .eret_d(eret_d), .n41364(n41364), .n41285(n41285), .load_d(load_d), 
            .n32910(n32910), .n32356(n32356), .n10(n10), .store_d(store_d), 
            .n41361(n41361), .break_d(break_d), .n41367(n41367), .valid_d(valid_d), 
            .n10_adj_145(n10_adj_6254), .n30070(n30070), .n41196(n41196), 
            .n30888(n30888), .n41291(n41291), .n41373(n41373), .n41208(n41208), 
            .n31207(n31207), .\instruction_d[13] (instruction_d[13]), .n31218(n31218), 
            .\instruction_d[12] (instruction_d[12]), .n31219(n31219), .n31542(n31542), 
            .branch_d(branch_d), .write_enable_d(write_enable_d), .n41227(n41227), 
            .n41229(n41229), .n41281(n41281), .\instruction_d[11] (instruction_d[11]), 
            .n31221(n31221), .n41377(n41377), .n31216(n31216), .n41376(n41376), 
            .n31212(n31212), .n41375(n41375), .n31220(n31220), .n31213(n31213), 
            .n41368(n41368), .n31217(n31217), .n41374(n41374), .n31214(n31214), 
            .n41371(n41371), .n31211(n31211), .n41372(n41372), .n31209(n31209), 
            .n41348(n41348), .n31206(n31206), .n41370(n41370), .n31210(n31210), 
            .n41369(n41369), .n31215(n31215), .\instruction_d[14] (instruction_d[14]), 
            .n31208(n31208), .branch_predict_taken_d(branch_predict_taken_d), 
            .n41179(n41179), .n30820(n30820), .n41175(n41175), .adder_op_d_N_1366(adder_op_d_N_1366), 
            .n6026(n6026), .n41187(n41187), .valid_f(valid_f), .n41203(n41203), 
            .n31132(n31132), .n45181(n45181), .valid_f_N_1250(valid_f_N_1250), 
            .bypass_data_1({bypass_data_1}), .n31309(n31309), .n31310(n31310), 
            .n31323(n31323), .n31298(n31298), .n31300(n31300), .n31322(n31322), 
            .n31302(n31302), .n31316(n31316), .n31304(n31304), .\extended_immediate[31] (extended_immediate[31]), 
            .n31320(n31320), .n31317(n31317), .n41452(n41452), .n31306(n31306), 
            .n31295(n31295), .n31311(n31311), .n31313(n31313), .n31315(n31315), 
            .n31319(n31319), .n31321(n31321), .n31296(n31296), .n31314(n31314), 
            .n31318(n31318), .n31308(n31308), .n31294(n31294), .n31325(n31325), 
            .n31312(n31312), .n31324(n31324), .n31297(n31297), .n31299(n31299), 
            .n31301(n31301), .n31303(n31303), .n31305(n31305), .n31307(n31307), 
            .x_bypass_enable_d(x_bypass_enable_d), .x_result_sel_csr_d(x_result_sel_csr_d), 
            .n41296(n41296), .n41248(n41248), .n41441(n41441), .n41319(n41319), 
            .n45105(n45105), .n41241(n41241), .n30216(n30216), .n31519(n31519), 
            .m_bypass_enable_d(m_bypass_enable_d), .n41408(n41408), .n6760(n6760), 
            .n2(n2_adj_6244), .n19987(n19987), .n31549(n31549), .n6761(n6761), 
            .n2_adj_146(n2_adj_6243), .n6762(n6762), .n2_adj_147(n2_adj_6242), 
            .n6763(n6763), .n2_adj_148(n2_adj_6241), .m_result_sel_compare_d(m_result_sel_compare_d), 
            .n41451(n41451), .n6768(n6768), .n6764(n6764), .n10589(n10589), 
            .n45183(n45183), .n40093(n40093), .n40094(n40094), .n6766(n6766), 
            .n10585(n10585), .n6769(n6769), .n10591(n10591), .n41419(n41419), 
            .n10485(n10485), .x_bypass_enable_x(x_bypass_enable_x), .n32006(n32006), 
            .m_bypass_enable_m(m_bypass_enable_m), .n31984(n31984), .n10593(n10593), 
            .n6767(n6767), .n10587(n10587), .n41312(n41312), .n41437(n41437), 
            .n41184(n41184), .n37939(n37939), .n41366(n41366), .n41201(n41201), 
            .\d_result_sel_1_d[1] (d_result_sel_1_d[1]), .n6771(n6771), 
            .n10595(n10595), .n37933(n37933), .n41205(n41205), .n37934(n37934), 
            .n37936(n37936), .n6765(n6765), .n10452(n10452), .n37937(n37937), 
            .n37938(n37938), .n37935(n37935), .n31494(n31494)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(899[14] 975[6])
    lm32_adder adder (.operand_0_x({operand_0_x}), .operand_1_x({operand_1_x[31:2], 
            \operand_1_x[1] , operand_1_x[0]}), .adder_op_x(adder_op_x), 
            .adder_op_x_n(adder_op_x_n), .adder_result_x({\adder_result_x[31] , 
            \adder_result_x[30] , \adder_result_x[29] , \adder_result_x[28] , 
            \adder_result_x[27] , \adder_result_x[26] , \adder_result_x[25] , 
            \adder_result_x[24] , \adder_result_x[23] , \adder_result_x[22] , 
            \adder_result_x[21] , \adder_result_x[20] , \adder_result_x[19] , 
            \adder_result_x[18] , \adder_result_x[17] , \adder_result_x[16] , 
            adder_result_x[15:0]}), .adder_carry_n_x(adder_carry_n_x)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1046[12] 1056[6])
    
endmodule
//
// Verilog Description of module lm32_shifter
//

module lm32_shifter (\operand_1_x[4] , \operand_1_x[3] , left_shift_result, 
            REF_CLK_c, REF_CLK_c_enable_1624, REF_CLK_c_enable_1606, \operand_1_x[2] , 
            \operand_1_x[1] , \operand_1_x[0] , operand_0_x, direction_x, 
            direction_m, \condition_x[2] , REF_CLK_c_enable_1030, \left_shift_result[27] , 
            \left_shift_result[25] , \left_shift_result[21] , \left_shift_result[10] , 
            \left_shift_result[6] , \left_shift_result[4] , \left_shift_result[0] , 
            \shifter_result_m[1] , \shifter_result_m[2] , \shifter_result_m[3] , 
            \shifter_result_m[5] , \shifter_result_m[7] , \shifter_result_m[8] , 
            \shifter_result_m[9] , \shifter_result_m[11] , \shifter_result_m[12] , 
            \shifter_result_m[13] , \shifter_result_m[14] , \shifter_result_m[15] , 
            \shifter_result_m[16] , \shifter_result_m[17] , \shifter_result_m[18] , 
            \shifter_result_m[19] , \shifter_result_m[20] , \shifter_result_m[22] , 
            \shifter_result_m[23] , \shifter_result_m[24] , \shifter_result_m[26] , 
            \shifter_result_m[28] , \shifter_result_m[29] , \shifter_result_m[30] ) /* synthesis syn_module_defined=1 */ ;
    input \operand_1_x[4] ;
    input \operand_1_x[3] ;
    output [31:0]left_shift_result;
    input REF_CLK_c;
    input REF_CLK_c_enable_1624;
    input REF_CLK_c_enable_1606;
    input \operand_1_x[2] ;
    input \operand_1_x[1] ;
    input \operand_1_x[0] ;
    input [31:0]operand_0_x;
    input direction_x;
    output direction_m;
    input \condition_x[2] ;
    input REF_CLK_c_enable_1030;
    output \left_shift_result[27] ;
    output \left_shift_result[25] ;
    output \left_shift_result[21] ;
    output \left_shift_result[10] ;
    output \left_shift_result[6] ;
    output \left_shift_result[4] ;
    output \left_shift_result[0] ;
    output \shifter_result_m[1] ;
    output \shifter_result_m[2] ;
    output \shifter_result_m[3] ;
    output \shifter_result_m[5] ;
    output \shifter_result_m[7] ;
    output \shifter_result_m[8] ;
    output \shifter_result_m[9] ;
    output \shifter_result_m[11] ;
    output \shifter_result_m[12] ;
    output \shifter_result_m[13] ;
    output \shifter_result_m[14] ;
    output \shifter_result_m[15] ;
    output \shifter_result_m[16] ;
    output \shifter_result_m[17] ;
    output \shifter_result_m[18] ;
    output \shifter_result_m[19] ;
    output \shifter_result_m[20] ;
    output \shifter_result_m[22] ;
    output \shifter_result_m[23] ;
    output \shifter_result_m[24] ;
    output \shifter_result_m[26] ;
    output \shifter_result_m[28] ;
    output \shifter_result_m[29] ;
    output \shifter_result_m[30] ;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    
    wire n208, n224;
    wire [63:0]left_shift_result_31__N_2627;
    
    wire n41063, n45195, n41060, n45197, n41053, n45198, n41048, 
        n45199, n41418, fill_value, n31, n223, n41404, n93, n94, 
        n207, n41043, n45200, n206, n222, n73, n77, n137, n81, 
        n85, n145, n41433;
    wire [31:0]right_shift_operand;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(96[23:42])
    
    wire n160, n9, n11, n6, n8, n70, n10, n12, n74, n78, 
        n138, n4, n5, n7, n69, n3, n72, n205, n221, n14, 
        n76, n71, n13, n75, n80, n140, n79, n139, n41678, 
        n89, n153, n36181, n36182, n152, n84, n144, n88, n92, 
        n24, n26, n28, n30, n16, n18, n20, n22;
    wire [31:0]left_shift_result_c;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(93[22:39])
    
    wire n146, n154, n41068, n41069, n41070, n156, n36062, n148, 
        n36061, n155, n36317, n147, n36316, n36053, n36052, n41072, 
        n41073, n41074, n41657, n45203, n41658, n45206, n45207, 
        n45208, n149, n157, n45209, n83, n143, n87, n91, n151, 
        n23, n25, n27, n29, n41679, n15, n17, n19, n21, n159, 
        n82, n142, n86, n90, n150, n32, n141, n41318, n41655, 
        n41656, n41271, n41327, n96, n41680, n158, n209, n210, 
        n211, n95, n212, n213, n214, n215, n216, n41042, n41059, 
        n41062, n41065, n41066;
    
    PFUMX shift_right_13_i272 (.BLUT(n208), .ALUT(n224), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2627[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;
    PFUMX i34304 (.BLUT(n41063), .ALUT(n45195), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2627[6]));
    PFUMX i34302 (.BLUT(n41060), .ALUT(n45197), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2627[7]));
    PFUMX i34300 (.BLUT(n41053), .ALUT(n45198), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2627[0]));
    PFUMX i34298 (.BLUT(n41048), .ALUT(n45199), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2627[1]));
    LUT4 i4178_3_lut_4_lut (.A(n41418), .B(\operand_1_x[3] ), .C(fill_value), 
         .D(n31), .Z(n223)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4178_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4192_3_lut_4_lut (.A(n41404), .B(\operand_1_x[4] ), .C(fill_value), 
         .D(n93), .Z(left_shift_result_31__N_2627[28])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4192_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4194_3_lut_4_lut (.A(n41404), .B(\operand_1_x[4] ), .C(fill_value), 
         .D(n94), .Z(left_shift_result_31__N_2627[29])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4194_3_lut_4_lut.init = 16'hf1e0;
    PFUMX shift_right_13_i271 (.BLUT(n207), .ALUT(n223), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2627[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;
    PFUMX i34296 (.BLUT(n41043), .ALUT(n45200), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2627[5]));
    FD1P3DX right_shift_result_i0_i0 (.D(left_shift_result_31__N_2627[0]), 
            .SP(REF_CLK_c_enable_1624), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i0.GSR = "ENABLED";
    PFUMX shift_right_13_i270 (.BLUT(n206), .ALUT(n222), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2627[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;
    LUT4 shift_right_13_i137_3_lut (.A(n73), .B(n77), .C(\operand_1_x[2] ), 
         .Z(n137)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i137_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i145_3_lut (.A(n81), .B(n85), .C(\operand_1_x[2] ), 
         .Z(n145)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i145_3_lut.init = 16'hcaca;
    LUT4 i4170_3_lut_4_lut (.A(n41433), .B(\operand_1_x[2] ), .C(fill_value), 
         .D(right_shift_operand[31]), .Z(n160)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4170_3_lut_4_lut.init = 16'hf1e0;
    LUT4 shift_right_13_i73_3_lut (.A(n9), .B(n11), .C(\operand_1_x[1] ), 
         .Z(n73)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i73_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i9_3_lut (.A(right_shift_operand[8]), .B(right_shift_operand[9]), 
         .C(\operand_1_x[0] ), .Z(n9)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i9_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i70_3_lut (.A(n6), .B(n8), .C(\operand_1_x[1] ), 
         .Z(n70)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i70_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i74_3_lut (.A(n10), .B(n12), .C(\operand_1_x[1] ), 
         .Z(n74)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i74_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i10_3_lut (.A(right_shift_operand[9]), .B(right_shift_operand[10]), 
         .C(\operand_1_x[0] ), .Z(n10)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i10_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i12_3_lut (.A(right_shift_operand[11]), .B(right_shift_operand[12]), 
         .C(\operand_1_x[0] ), .Z(n12)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i12_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i6_3_lut (.A(right_shift_operand[5]), .B(right_shift_operand[6]), 
         .C(\operand_1_x[0] ), .Z(n6)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i6_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i8_3_lut (.A(right_shift_operand[7]), .B(right_shift_operand[8]), 
         .C(\operand_1_x[0] ), .Z(n8)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i8_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i6_3_lut (.A(operand_0_x[5]), .B(operand_0_x[26]), 
         .C(direction_x), .Z(right_shift_operand[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i6_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i7_3_lut (.A(operand_0_x[6]), .B(operand_0_x[25]), 
         .C(direction_x), .Z(right_shift_operand[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i7_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i8_3_lut (.A(operand_0_x[7]), .B(operand_0_x[24]), 
         .C(direction_x), .Z(right_shift_operand[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i8_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i138_3_lut (.A(n74), .B(n78), .C(\operand_1_x[2] ), 
         .Z(n138)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i138_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i4_3_lut (.A(right_shift_operand[3]), .B(right_shift_operand[4]), 
         .C(\operand_1_x[0] ), .Z(n4)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i4_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i4_3_lut (.A(operand_0_x[3]), .B(operand_0_x[28]), 
         .C(direction_x), .Z(right_shift_operand[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i4_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i5_3_lut (.A(operand_0_x[4]), .B(operand_0_x[27]), 
         .C(direction_x), .Z(right_shift_operand[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i5_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i2_3_lut (.A(operand_0_x[1]), .B(operand_0_x[30]), 
         .C(direction_x), .Z(right_shift_operand[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i2_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i3_3_lut (.A(operand_0_x[2]), .B(operand_0_x[29]), 
         .C(direction_x), .Z(right_shift_operand[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i3_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i69_3_lut (.A(n5), .B(n7), .C(\operand_1_x[1] ), 
         .Z(n69)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i69_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i3_3_lut (.A(right_shift_operand[2]), .B(right_shift_operand[3]), 
         .C(\operand_1_x[0] ), .Z(n3)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i3_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i5_3_lut (.A(right_shift_operand[4]), .B(right_shift_operand[5]), 
         .C(\operand_1_x[0] ), .Z(n5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i5_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i7_3_lut (.A(right_shift_operand[6]), .B(right_shift_operand[7]), 
         .C(\operand_1_x[0] ), .Z(n7)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i7_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i11_3_lut (.A(right_shift_operand[10]), .B(right_shift_operand[11]), 
         .C(\operand_1_x[0] ), .Z(n11)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i11_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i9_3_lut (.A(operand_0_x[8]), .B(operand_0_x[23]), 
         .C(direction_x), .Z(right_shift_operand[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i9_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i72_3_lut (.A(n8), .B(n10), .C(\operand_1_x[1] ), 
         .Z(n72)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i72_3_lut.init = 16'hcaca;
    PFUMX shift_right_13_i269 (.BLUT(n205), .ALUT(n221), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2627[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;
    LUT4 shift_right_13_i76_3_lut (.A(n12), .B(n14), .C(\operand_1_x[1] ), 
         .Z(n76)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i76_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i71_3_lut (.A(n7), .B(n9), .C(\operand_1_x[1] ), 
         .Z(n71)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i71_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i75_3_lut (.A(n11), .B(n13), .C(\operand_1_x[1] ), 
         .Z(n75)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i75_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i140_3_lut (.A(n76), .B(n80), .C(\operand_1_x[2] ), 
         .Z(n140)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i140_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i139_3_lut (.A(n75), .B(n79), .C(\operand_1_x[2] ), 
         .Z(n139)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i139_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i10_3_lut (.A(operand_0_x[9]), .B(operand_0_x[22]), 
         .C(direction_x), .Z(right_shift_operand[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i10_3_lut.init = 16'hcaca;
    LUT4 n4_bdd_3_lut (.A(right_shift_operand[2]), .B(right_shift_operand[1]), 
         .C(\operand_1_x[0] ), .Z(n41678)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n4_bdd_3_lut.init = 16'hacac;
    LUT4 operand_0_x_31__I_0_22_i11_3_lut (.A(operand_0_x[10]), .B(operand_0_x[21]), 
         .C(direction_x), .Z(right_shift_operand[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i11_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i12_3_lut (.A(operand_0_x[11]), .B(operand_0_x[20]), 
         .C(direction_x), .Z(right_shift_operand[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i12_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i153_3_lut (.A(n89), .B(n93), .C(\operand_1_x[2] ), 
         .Z(n153)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i153_3_lut.init = 16'hcaca;
    PFUMX i31011 (.BLUT(n36181), .ALUT(n36182), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2627[8]));
    FD1P3DX direction_m_20 (.D(direction_x), .SP(REF_CLK_c_enable_1624), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(direction_m)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam direction_m_20.GSR = "ENABLED";
    LUT4 shift_right_13_i216_3_lut_rep_1152 (.A(n152), .B(n160), .C(\operand_1_x[3] ), 
         .Z(n45197)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i216_3_lut_rep_1152.init = 16'hcaca;
    LUT4 shift_right_13_i209_3_lut_rep_1153 (.A(n145), .B(n153), .C(\operand_1_x[3] ), 
         .Z(n45198)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i209_3_lut_rep_1153.init = 16'hcaca;
    LUT4 shift_right_13_i144_3_lut (.A(n80), .B(n84), .C(\operand_1_x[2] ), 
         .Z(n144)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i144_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i152_3_lut (.A(n88), .B(n92), .C(\operand_1_x[2] ), 
         .Z(n152)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i152_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i88_3_lut (.A(n24), .B(n26), .C(\operand_1_x[1] ), 
         .Z(n88)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i88_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i92_3_lut (.A(n28), .B(n30), .C(\operand_1_x[1] ), 
         .Z(n92)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i92_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i28_3_lut (.A(right_shift_operand[27]), .B(right_shift_operand[28]), 
         .C(\operand_1_x[0] ), .Z(n28)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i28_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i30_3_lut (.A(right_shift_operand[29]), .B(right_shift_operand[30]), 
         .C(\operand_1_x[0] ), .Z(n30)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i30_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i30_3_lut (.A(operand_0_x[29]), .B(operand_0_x[2]), 
         .C(direction_x), .Z(right_shift_operand[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i30_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i31_3_lut (.A(operand_0_x[30]), .B(operand_0_x[1]), 
         .C(direction_x), .Z(right_shift_operand[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i31_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i28_3_lut (.A(operand_0_x[27]), .B(operand_0_x[4]), 
         .C(direction_x), .Z(right_shift_operand[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i28_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i29_3_lut (.A(operand_0_x[28]), .B(operand_0_x[3]), 
         .C(direction_x), .Z(right_shift_operand[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i29_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i80_3_lut (.A(n16), .B(n18), .C(\operand_1_x[1] ), 
         .Z(n80)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i80_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i84_3_lut (.A(n20), .B(n22), .C(\operand_1_x[1] ), 
         .Z(n84)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i84_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i20_3_lut (.A(right_shift_operand[19]), .B(right_shift_operand[20]), 
         .C(\operand_1_x[0] ), .Z(n20)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i20_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i22_3_lut (.A(right_shift_operand[21]), .B(right_shift_operand[22]), 
         .C(\operand_1_x[0] ), .Z(n22)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i22_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i16_4_lut (.A(operand_0_x[15]), .B(operand_0_x[16]), 
         .C(direction_x), .D(\operand_1_x[0] ), .Z(n16)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A !((C (D)+!C !(D))+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i16_4_lut.init = 16'hacca;
    LUT4 shift_right_13_i18_3_lut (.A(right_shift_operand[17]), .B(right_shift_operand[18]), 
         .C(\operand_1_x[0] ), .Z(n18)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i18_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i18_3_lut (.A(operand_0_x[17]), .B(operand_0_x[14]), 
         .C(direction_x), .Z(right_shift_operand[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i18_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i19_3_lut (.A(operand_0_x[18]), .B(operand_0_x[13]), 
         .C(direction_x), .Z(right_shift_operand[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i19_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i22_3_lut (.A(operand_0_x[21]), .B(operand_0_x[10]), 
         .C(direction_x), .Z(right_shift_operand[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i22_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i23_3_lut (.A(operand_0_x[22]), .B(operand_0_x[9]), 
         .C(direction_x), .Z(right_shift_operand[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i23_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i20_3_lut (.A(operand_0_x[19]), .B(operand_0_x[12]), 
         .C(direction_x), .Z(right_shift_operand[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i20_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i21_3_lut (.A(operand_0_x[20]), .B(operand_0_x[11]), 
         .C(direction_x), .Z(right_shift_operand[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i21_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i24_3_lut (.A(right_shift_operand[23]), .B(right_shift_operand[24]), 
         .C(\operand_1_x[0] ), .Z(n24)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i24_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i26_3_lut (.A(right_shift_operand[25]), .B(right_shift_operand[26]), 
         .C(\operand_1_x[0] ), .Z(n26)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i26_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i26_3_lut (.A(operand_0_x[25]), .B(operand_0_x[6]), 
         .C(direction_x), .Z(right_shift_operand[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i26_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i27_3_lut (.A(operand_0_x[26]), .B(operand_0_x[5]), 
         .C(direction_x), .Z(right_shift_operand[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i27_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i24_3_lut (.A(operand_0_x[23]), .B(operand_0_x[8]), 
         .C(direction_x), .Z(right_shift_operand[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i24_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i25_3_lut (.A(operand_0_x[24]), .B(operand_0_x[7]), 
         .C(direction_x), .Z(right_shift_operand[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i25_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i32_3_lut (.A(operand_0_x[31]), .B(operand_0_x[0]), 
         .C(direction_x), .Z(right_shift_operand[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i32_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[31]), 
         .Z(fill_value)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(116[21] 118[29])
    defparam i1_3_lut.init = 16'h2020;
    FD1P3DX right_shift_result_i0_i1 (.D(left_shift_result_31__N_2627[1]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i1.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i2 (.D(left_shift_result_31__N_2627[2]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i2.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i3 (.D(left_shift_result_31__N_2627[3]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i3.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i4 (.D(left_shift_result_31__N_2627[4]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\left_shift_result[27] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i4.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i5 (.D(left_shift_result_31__N_2627[5]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i5.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i6 (.D(left_shift_result_31__N_2627[6]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\left_shift_result[25] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i6.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i7 (.D(left_shift_result_31__N_2627[7]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i7.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i8 (.D(left_shift_result_31__N_2627[8]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i8.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i9 (.D(left_shift_result_31__N_2627[9]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i9.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i10 (.D(left_shift_result_31__N_2627[10]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\left_shift_result[21] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i10.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i11 (.D(left_shift_result_31__N_2627[11]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i11.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i12 (.D(left_shift_result_31__N_2627[12]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i12.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i13 (.D(left_shift_result_31__N_2627[13]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i13.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i14 (.D(left_shift_result_31__N_2627[14]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i14.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i15 (.D(left_shift_result_31__N_2627[15]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i15.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i16 (.D(left_shift_result_31__N_2627[16]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i16.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i17 (.D(left_shift_result_31__N_2627[17]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i17.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i18 (.D(left_shift_result_31__N_2627[18]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i18.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i19 (.D(left_shift_result_31__N_2627[19]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i19.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i20 (.D(left_shift_result_31__N_2627[20]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i20.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i21 (.D(left_shift_result_31__N_2627[21]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\left_shift_result[10] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i21.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i22 (.D(left_shift_result_31__N_2627[22]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i22.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i23 (.D(left_shift_result_31__N_2627[23]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i23.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i24 (.D(left_shift_result_31__N_2627[24]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i24.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i25 (.D(left_shift_result_31__N_2627[25]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\left_shift_result[6] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i25.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i26 (.D(left_shift_result_31__N_2627[26]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i26.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i27 (.D(left_shift_result_31__N_2627[27]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\left_shift_result[4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i27.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i28 (.D(left_shift_result_31__N_2627[28]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i28.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i29 (.D(left_shift_result_31__N_2627[29]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i29.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i30 (.D(left_shift_result_31__N_2627[30]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(left_shift_result_c[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i30.GSR = "ENABLED";
    FD1P3DX right_shift_result_i0_i31 (.D(left_shift_result_31__N_2627[31]), 
            .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\left_shift_result[0] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i31.GSR = "ENABLED";
    LUT4 shift_right_13_i210_3_lut_rep_1154 (.A(n146), .B(n154), .C(\operand_1_x[3] ), 
         .Z(n45199)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i210_3_lut_rep_1154.init = 16'hcaca;
    LUT4 n72_bdd_3_lut_35839 (.A(n4), .B(n6), .C(\operand_1_x[1] ), .Z(n41068)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n72_bdd_3_lut_35839.init = 16'hcaca;
    LUT4 n41068_bdd_3_lut (.A(n41068), .B(n72), .C(\operand_1_x[2] ), 
         .Z(n41069)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41068_bdd_3_lut.init = 16'hcaca;
    LUT4 n41069_bdd_3_lut (.A(n41069), .B(n140), .C(\operand_1_x[3] ), 
         .Z(n41070)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41069_bdd_3_lut.init = 16'hcaca;
    LUT4 i30890_3_lut (.A(n156), .B(fill_value), .C(\operand_1_x[3] ), 
         .Z(n36062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30890_3_lut.init = 16'hcaca;
    LUT4 i30889_3_lut (.A(n140), .B(n148), .C(\operand_1_x[3] ), .Z(n36061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30889_3_lut.init = 16'hcaca;
    LUT4 i31145_3_lut (.A(n155), .B(fill_value), .C(\operand_1_x[3] ), 
         .Z(n36317)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31145_3_lut.init = 16'hcaca;
    LUT4 i31144_3_lut (.A(n139), .B(n147), .C(\operand_1_x[3] ), .Z(n36316)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31144_3_lut.init = 16'hcaca;
    LUT4 i30881_3_lut (.A(n154), .B(fill_value), .C(\operand_1_x[3] ), 
         .Z(n36053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30881_3_lut.init = 16'hcaca;
    LUT4 i30880_3_lut (.A(n138), .B(n146), .C(\operand_1_x[3] ), .Z(n36052)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30880_3_lut.init = 16'hcaca;
    LUT4 n71_bdd_3_lut_35759 (.A(n3), .B(n5), .C(\operand_1_x[1] ), .Z(n41072)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n71_bdd_3_lut_35759.init = 16'hcaca;
    LUT4 n41072_bdd_3_lut (.A(n41072), .B(n71), .C(\operand_1_x[2] ), 
         .Z(n41073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41072_bdd_3_lut.init = 16'hcaca;
    LUT4 n41073_bdd_3_lut (.A(n41073), .B(n139), .C(\operand_1_x[3] ), 
         .Z(n41074)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41073_bdd_3_lut.init = 16'hcaca;
    PFUMX i34469 (.BLUT(n41657), .ALUT(n45203), .C0(\operand_1_x[2] ), 
          .Z(n41658));
    LUT4 shift_right_13_i69_3_lut_rep_1158 (.A(n5), .B(n7), .C(\operand_1_x[1] ), 
         .Z(n45203)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i69_3_lut_rep_1158.init = 16'hcaca;
    LUT4 shift_right_13_i70_3_lut_rep_1161 (.A(n6), .B(n8), .C(\operand_1_x[1] ), 
         .Z(n45206)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i70_3_lut_rep_1161.init = 16'hcaca;
    LUT4 shift_right_13_i211_3_lut_rep_1162 (.A(n147), .B(n155), .C(\operand_1_x[3] ), 
         .Z(n45207)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i211_3_lut_rep_1162.init = 16'hcaca;
    LUT4 shift_right_13_i212_3_lut_rep_1163 (.A(n148), .B(n156), .C(\operand_1_x[3] ), 
         .Z(n45208)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i212_3_lut_rep_1163.init = 16'hcaca;
    LUT4 shift_right_13_i213_3_lut_rep_1164 (.A(n149), .B(n157), .C(\operand_1_x[3] ), 
         .Z(n45209)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i213_3_lut_rep_1164.init = 16'hcaca;
    LUT4 shift_right_13_i143_3_lut (.A(n79), .B(n83), .C(\operand_1_x[2] ), 
         .Z(n143)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i143_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i151_3_lut (.A(n87), .B(n91), .C(\operand_1_x[2] ), 
         .Z(n151)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i151_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i87_3_lut (.A(n23), .B(n25), .C(\operand_1_x[1] ), 
         .Z(n87)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i87_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i91_3_lut (.A(n27), .B(n29), .C(\operand_1_x[1] ), 
         .Z(n91)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i91_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i27_3_lut (.A(right_shift_operand[26]), .B(right_shift_operand[27]), 
         .C(\operand_1_x[0] ), .Z(n27)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i27_3_lut.init = 16'hcaca;
    LUT4 n41678_bdd_3_lut (.A(n41678), .B(n4), .C(\operand_1_x[1] ), .Z(n41679)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41678_bdd_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i29_3_lut (.A(right_shift_operand[28]), .B(right_shift_operand[29]), 
         .C(\operand_1_x[0] ), .Z(n29)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i29_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i79_3_lut (.A(n15), .B(n17), .C(\operand_1_x[1] ), 
         .Z(n79)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i79_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i83_3_lut (.A(n19), .B(n21), .C(\operand_1_x[1] ), 
         .Z(n83)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i83_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i19_3_lut (.A(right_shift_operand[18]), .B(right_shift_operand[19]), 
         .C(\operand_1_x[0] ), .Z(n19)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i19_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i21_3_lut (.A(right_shift_operand[20]), .B(right_shift_operand[21]), 
         .C(\operand_1_x[0] ), .Z(n21)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i21_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i15_3_lut (.A(right_shift_operand[14]), .B(right_shift_operand[15]), 
         .C(\operand_1_x[0] ), .Z(n15)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i15_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i16_3_lut (.A(operand_0_x[15]), .B(operand_0_x[16]), 
         .C(direction_x), .Z(right_shift_operand[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i16_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i17_3_lut (.A(right_shift_operand[16]), .B(right_shift_operand[17]), 
         .C(\operand_1_x[0] ), .Z(n17)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i17_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i17_3_lut (.A(operand_0_x[16]), .B(operand_0_x[15]), 
         .C(direction_x), .Z(right_shift_operand[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i17_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i15_3_lut (.A(operand_0_x[14]), .B(operand_0_x[17]), 
         .C(direction_x), .Z(right_shift_operand[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i15_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i23_3_lut (.A(right_shift_operand[22]), .B(right_shift_operand[23]), 
         .C(\operand_1_x[0] ), .Z(n23)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i23_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i25_3_lut (.A(right_shift_operand[24]), .B(right_shift_operand[25]), 
         .C(\operand_1_x[0] ), .Z(n25)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i25_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i31_3_lut (.A(right_shift_operand[30]), .B(right_shift_operand[31]), 
         .C(\operand_1_x[0] ), .Z(n31)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i31_3_lut.init = 16'hcaca;
    LUT4 i4184_3_lut_4_lut (.A(\operand_1_x[3] ), .B(\operand_1_x[4] ), 
         .C(fill_value), .D(n153), .Z(left_shift_result_31__N_2627[24])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4184_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4186_3_lut_4_lut (.A(\operand_1_x[3] ), .B(\operand_1_x[4] ), 
         .C(fill_value), .D(n154), .Z(left_shift_result_31__N_2627[25])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4186_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4188_3_lut_4_lut (.A(\operand_1_x[3] ), .B(\operand_1_x[4] ), 
         .C(fill_value), .D(n155), .Z(left_shift_result_31__N_2627[26])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4188_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4190_3_lut_4_lut (.A(\operand_1_x[3] ), .B(\operand_1_x[4] ), 
         .C(fill_value), .D(n156), .Z(left_shift_result_31__N_2627[27])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4190_3_lut_4_lut.init = 16'hf1e0;
    LUT4 shift_right_13_i215_3_lut_rep_1150 (.A(n151), .B(n159), .C(\operand_1_x[3] ), 
         .Z(n45195)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i215_3_lut_rep_1150.init = 16'hcaca;
    LUT4 shift_right_13_i142_3_lut (.A(n78), .B(n82), .C(\operand_1_x[2] ), 
         .Z(n142)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i142_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i150_3_lut (.A(n86), .B(n90), .C(\operand_1_x[2] ), 
         .Z(n150)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i150_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i86_3_lut (.A(n22), .B(n24), .C(\operand_1_x[1] ), 
         .Z(n86)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i86_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i90_3_lut (.A(n26), .B(n28), .C(\operand_1_x[1] ), 
         .Z(n90)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i90_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i78_3_lut (.A(n14), .B(n16), .C(\operand_1_x[1] ), 
         .Z(n78)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i78_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i82_3_lut (.A(n18), .B(n20), .C(\operand_1_x[1] ), 
         .Z(n82)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i82_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i14_3_lut (.A(right_shift_operand[13]), .B(right_shift_operand[14]), 
         .C(\operand_1_x[0] ), .Z(n14)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i14_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i14_3_lut (.A(operand_0_x[13]), .B(operand_0_x[18]), 
         .C(direction_x), .Z(right_shift_operand[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i14_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i94_3_lut (.A(n30), .B(n32), .C(\operand_1_x[1] ), 
         .Z(n94)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i94_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i32_3_lut (.A(right_shift_operand[31]), .B(fill_value), 
         .C(\operand_1_x[0] ), .Z(n32)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i32_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i141_3_lut (.A(n77), .B(n81), .C(\operand_1_x[2] ), 
         .Z(n141)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i141_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i149_3_lut (.A(n85), .B(n89), .C(\operand_1_x[2] ), 
         .Z(n149)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i149_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i85_3_lut (.A(n21), .B(n23), .C(\operand_1_x[1] ), 
         .Z(n85)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i85_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i89_3_lut (.A(n25), .B(n27), .C(\operand_1_x[1] ), 
         .Z(n89)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i89_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i77_3_lut (.A(n13), .B(n15), .C(\operand_1_x[1] ), 
         .Z(n77)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i77_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i81_3_lut (.A(n17), .B(n19), .C(\operand_1_x[1] ), 
         .Z(n81)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i81_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i13_3_lut (.A(right_shift_operand[12]), .B(right_shift_operand[13]), 
         .C(\operand_1_x[0] ), .Z(n13)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i13_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i13_3_lut (.A(operand_0_x[12]), .B(operand_0_x[19]), 
         .C(direction_x), .Z(right_shift_operand[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i13_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i93_3_lut (.A(n29), .B(n31), .C(\operand_1_x[1] ), 
         .Z(n93)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i93_3_lut.init = 16'hcaca;
    LUT4 i4173_2_lut_rep_999 (.A(\operand_1_x[2] ), .B(\operand_1_x[3] ), 
         .Z(n41404)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4173_2_lut_rep_999.init = 16'heeee;
    LUT4 i4174_3_lut_4_lut (.A(\operand_1_x[2] ), .B(\operand_1_x[3] ), 
         .C(fill_value), .D(n93), .Z(n221)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4174_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4176_3_lut_4_lut (.A(\operand_1_x[2] ), .B(\operand_1_x[3] ), 
         .C(fill_value), .D(n94), .Z(n222)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4176_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4167_2_lut_rep_1013 (.A(\operand_1_x[1] ), .B(\operand_1_x[2] ), 
         .Z(n41418)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4167_2_lut_rep_1013.init = 16'heeee;
    LUT4 i4177_2_lut_rep_913_3_lut (.A(\operand_1_x[1] ), .B(\operand_1_x[2] ), 
         .C(\operand_1_x[3] ), .Z(n41318)) /* synthesis lut_function=(A+(B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4177_2_lut_rep_913_3_lut.init = 16'hfefe;
    LUT4 i4168_3_lut_4_lut (.A(\operand_1_x[1] ), .B(\operand_1_x[2] ), 
         .C(fill_value), .D(n31), .Z(n159)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4168_3_lut_4_lut.init = 16'hf1e0;
    LUT4 right_shift_operand_1__bdd_3_lut_34482 (.A(operand_0_x[31]), .B(operand_0_x[0]), 
         .C(direction_x), .Z(n41655)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam right_shift_operand_1__bdd_3_lut_34482.init = 16'hacac;
    LUT4 n41655_bdd_3_lut (.A(n41655), .B(right_shift_operand[1]), .C(\operand_1_x[0] ), 
         .Z(n41656)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41655_bdd_3_lut.init = 16'hcaca;
    LUT4 n41656_bdd_3_lut (.A(n41656), .B(n3), .C(\operand_1_x[1] ), .Z(n41657)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41656_bdd_3_lut.init = 16'hcaca;
    LUT4 i4164_2_lut_rep_1028 (.A(\operand_1_x[0] ), .B(\operand_1_x[1] ), 
         .Z(n41433)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4164_2_lut_rep_1028.init = 16'heeee;
    LUT4 i4179_2_lut_rep_866_3_lut_4_lut (.A(\operand_1_x[0] ), .B(\operand_1_x[1] ), 
         .C(\operand_1_x[3] ), .D(\operand_1_x[2] ), .Z(n41271)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4179_2_lut_rep_866_3_lut_4_lut.init = 16'hfffe;
    LUT4 i4169_2_lut_rep_922_3_lut (.A(\operand_1_x[0] ), .B(\operand_1_x[1] ), 
         .C(\operand_1_x[2] ), .Z(n41327)) /* synthesis lut_function=(A+(B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4169_2_lut_rep_922_3_lut.init = 16'hfefe;
    LUT4 i4165_3_lut_4_lut (.A(\operand_1_x[0] ), .B(\operand_1_x[1] ), 
         .C(fill_value), .D(right_shift_operand[31]), .Z(n96)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4165_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i34486 (.BLUT(n41679), .ALUT(n45206), .C0(\operand_1_x[2] ), 
          .Z(n41680));
    LUT4 i31010_3_lut (.A(n153), .B(fill_value), .C(\operand_1_x[3] ), 
         .Z(n36182)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31010_3_lut.init = 16'hcaca;
    LUT4 i31009_3_lut (.A(n137), .B(n145), .C(\operand_1_x[3] ), .Z(n36181)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31009_3_lut.init = 16'hcaca;
    LUT4 i4180_3_lut_4_lut (.A(n41327), .B(\operand_1_x[3] ), .C(fill_value), 
         .D(right_shift_operand[31]), .Z(n224)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4180_3_lut_4_lut.init = 16'hf1e0;
    LUT4 left_shift_result_0__I_0_21_i2_3_lut (.A(left_shift_result_c[30]), 
         .B(left_shift_result_c[1]), .C(direction_m), .Z(\shifter_result_m[1] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i2_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i3_3_lut (.A(left_shift_result_c[29]), 
         .B(left_shift_result_c[2]), .C(direction_m), .Z(\shifter_result_m[2] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i3_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i4_3_lut (.A(left_shift_result_c[28]), 
         .B(left_shift_result_c[3]), .C(direction_m), .Z(\shifter_result_m[3] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i4_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i6_3_lut (.A(left_shift_result_c[26]), 
         .B(left_shift_result_c[5]), .C(direction_m), .Z(\shifter_result_m[5] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i6_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i8_3_lut (.A(left_shift_result_c[24]), 
         .B(left_shift_result_c[7]), .C(direction_m), .Z(\shifter_result_m[7] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i8_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i9_3_lut (.A(left_shift_result_c[23]), 
         .B(left_shift_result_c[8]), .C(direction_m), .Z(\shifter_result_m[8] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i9_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i10_3_lut (.A(left_shift_result_c[22]), 
         .B(left_shift_result_c[9]), .C(direction_m), .Z(\shifter_result_m[9] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i10_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i12_3_lut (.A(left_shift_result_c[20]), 
         .B(left_shift_result_c[11]), .C(direction_m), .Z(\shifter_result_m[11] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i12_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i13_3_lut (.A(left_shift_result_c[19]), 
         .B(left_shift_result_c[12]), .C(direction_m), .Z(\shifter_result_m[12] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i13_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i14_3_lut (.A(left_shift_result_c[18]), 
         .B(left_shift_result_c[13]), .C(direction_m), .Z(\shifter_result_m[13] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i14_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i15_3_lut (.A(left_shift_result_c[17]), 
         .B(left_shift_result_c[14]), .C(direction_m), .Z(\shifter_result_m[14] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i15_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i16_3_lut (.A(left_shift_result_c[16]), 
         .B(left_shift_result_c[15]), .C(direction_m), .Z(\shifter_result_m[15] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i16_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i17_3_lut (.A(left_shift_result_c[15]), 
         .B(left_shift_result_c[16]), .C(direction_m), .Z(\shifter_result_m[16] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i17_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i18_3_lut (.A(left_shift_result_c[14]), 
         .B(left_shift_result_c[17]), .C(direction_m), .Z(\shifter_result_m[17] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i18_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i19_3_lut (.A(left_shift_result_c[13]), 
         .B(left_shift_result_c[18]), .C(direction_m), .Z(\shifter_result_m[18] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i19_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i20_3_lut (.A(left_shift_result_c[12]), 
         .B(left_shift_result_c[19]), .C(direction_m), .Z(\shifter_result_m[19] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i20_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i21_3_lut (.A(left_shift_result_c[11]), 
         .B(left_shift_result_c[20]), .C(direction_m), .Z(\shifter_result_m[20] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i21_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i23_3_lut (.A(left_shift_result_c[9]), 
         .B(left_shift_result_c[22]), .C(direction_m), .Z(\shifter_result_m[22] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i23_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i24_3_lut (.A(left_shift_result_c[8]), 
         .B(left_shift_result_c[23]), .C(direction_m), .Z(\shifter_result_m[23] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i24_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i25_3_lut (.A(left_shift_result_c[7]), 
         .B(left_shift_result_c[24]), .C(direction_m), .Z(\shifter_result_m[24] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i25_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i205_3_lut (.A(n141), .B(n149), .C(\operand_1_x[3] ), 
         .Z(n205)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i205_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i27_3_lut (.A(left_shift_result_c[5]), 
         .B(left_shift_result_c[26]), .C(direction_m), .Z(\shifter_result_m[26] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i27_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i29_3_lut (.A(left_shift_result_c[3]), 
         .B(left_shift_result_c[28]), .C(direction_m), .Z(\shifter_result_m[28] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i29_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i30_3_lut (.A(left_shift_result_c[2]), 
         .B(left_shift_result_c[29]), .C(direction_m), .Z(\shifter_result_m[29] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i30_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i31_3_lut (.A(left_shift_result_c[1]), 
         .B(left_shift_result_c[30]), .C(direction_m), .Z(\shifter_result_m[30] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i31_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i214_3_lut_rep_1155 (.A(n150), .B(n158), .C(\operand_1_x[3] ), 
         .Z(n45200)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i214_3_lut_rep_1155.init = 16'hcaca;
    LUT4 shift_right_13_i206_3_lut (.A(n142), .B(n150), .C(\operand_1_x[3] ), 
         .Z(n206)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i206_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i273_3_lut (.A(n209), .B(fill_value), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2627[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i273_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i209_3_lut (.A(n145), .B(n153), .C(\operand_1_x[3] ), 
         .Z(n209)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i209_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i274_3_lut (.A(n210), .B(fill_value), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2627[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i274_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i210_3_lut (.A(n146), .B(n154), .C(\operand_1_x[3] ), 
         .Z(n210)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i210_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i146_3_lut (.A(n82), .B(n86), .C(\operand_1_x[2] ), 
         .Z(n146)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i146_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i154_3_lut (.A(n90), .B(n94), .C(\operand_1_x[2] ), 
         .Z(n154)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i154_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i275_3_lut (.A(n211), .B(fill_value), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2627[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i275_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i211_3_lut (.A(n147), .B(n155), .C(\operand_1_x[3] ), 
         .Z(n211)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i211_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i147_3_lut (.A(n83), .B(n87), .C(\operand_1_x[2] ), 
         .Z(n147)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i147_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i155_3_lut (.A(n91), .B(n95), .C(\operand_1_x[2] ), 
         .Z(n155)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i155_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i95_3_lut (.A(n31), .B(fill_value), .C(\operand_1_x[1] ), 
         .Z(n95)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i95_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i276_3_lut (.A(n212), .B(fill_value), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2627[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i276_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i212_3_lut (.A(n148), .B(n156), .C(\operand_1_x[3] ), 
         .Z(n212)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i212_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i148_3_lut (.A(n84), .B(n88), .C(\operand_1_x[2] ), 
         .Z(n148)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i148_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i156_3_lut (.A(n92), .B(n96), .C(\operand_1_x[2] ), 
         .Z(n156)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i156_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i277_3_lut (.A(n213), .B(fill_value), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2627[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i277_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i213_3_lut (.A(n149), .B(n157), .C(\operand_1_x[3] ), 
         .Z(n213)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i213_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i157_3_lut (.A(n93), .B(fill_value), .C(\operand_1_x[2] ), 
         .Z(n157)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i157_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i278_3_lut (.A(n214), .B(fill_value), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2627[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i278_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i214_3_lut (.A(n150), .B(n158), .C(\operand_1_x[3] ), 
         .Z(n214)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i214_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i158_3_lut (.A(n94), .B(fill_value), .C(\operand_1_x[2] ), 
         .Z(n158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i158_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i279_3_lut (.A(n215), .B(fill_value), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2627[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i279_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i215_3_lut (.A(n151), .B(n159), .C(\operand_1_x[3] ), 
         .Z(n215)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i215_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i280_3_lut (.A(n216), .B(fill_value), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2627[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i280_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i216_3_lut (.A(n152), .B(n160), .C(\operand_1_x[3] ), 
         .Z(n216)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i216_3_lut.init = 16'hcaca;
    LUT4 i4196_4_lut (.A(n31), .B(fill_value), .C(n41318), .D(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2627[30])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4196_4_lut.init = 16'hccca;
    LUT4 i4198_4_lut (.A(right_shift_operand[31]), .B(fill_value), .C(n41271), 
         .D(\operand_1_x[4] ), .Z(left_shift_result_31__N_2627[31])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i4198_4_lut.init = 16'hccca;
    LUT4 n41042_bdd_3_lut (.A(n41042), .B(n142), .C(\operand_1_x[3] ), 
         .Z(n41043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41042_bdd_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i207_3_lut (.A(n143), .B(n151), .C(\operand_1_x[3] ), 
         .Z(n207)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i207_3_lut.init = 16'hcaca;
    LUT4 n142_bdd_3_lut (.A(n70), .B(n74), .C(\operand_1_x[2] ), .Z(n41042)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n142_bdd_3_lut.init = 16'hcaca;
    LUT4 n41047_bdd_3_lut (.A(n41680), .B(n138), .C(\operand_1_x[3] ), 
         .Z(n41048)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41047_bdd_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i208_3_lut (.A(n144), .B(n152), .C(\operand_1_x[3] ), 
         .Z(n208)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i208_3_lut.init = 16'hcaca;
    LUT4 n41052_bdd_3_lut (.A(n41658), .B(n137), .C(\operand_1_x[3] ), 
         .Z(n41053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41052_bdd_3_lut.init = 16'hcaca;
    LUT4 n41059_bdd_3_lut (.A(n41059), .B(n144), .C(\operand_1_x[3] ), 
         .Z(n41060)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41059_bdd_3_lut.init = 16'hcaca;
    LUT4 n144_bdd_3_lut_34452 (.A(n72), .B(n76), .C(\operand_1_x[2] ), 
         .Z(n41059)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n144_bdd_3_lut_34452.init = 16'hcaca;
    LUT4 n143_bdd_3_lut_34500 (.A(n71), .B(n75), .C(\operand_1_x[2] ), 
         .Z(n41062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n143_bdd_3_lut_34500.init = 16'hcaca;
    LUT4 n41062_bdd_3_lut (.A(n41062), .B(n143), .C(\operand_1_x[3] ), 
         .Z(n41063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41062_bdd_3_lut.init = 16'hcaca;
    LUT4 n141_bdd_3_lut (.A(n69), .B(n73), .C(\operand_1_x[2] ), .Z(n41065)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n141_bdd_3_lut.init = 16'hcaca;
    LUT4 n41065_bdd_3_lut (.A(n41065), .B(n141), .C(\operand_1_x[3] ), 
         .Z(n41066)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41065_bdd_3_lut.init = 16'hcaca;
    PFUMX i34310 (.BLUT(n41074), .ALUT(n45207), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2627[2]));
    PFUMX i34308 (.BLUT(n41070), .ALUT(n45208), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2627[3]));
    PFUMX i30882 (.BLUT(n36052), .ALUT(n36053), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2627[9]));
    PFUMX i31146 (.BLUT(n36316), .ALUT(n36317), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2627[10]));
    PFUMX i30891 (.BLUT(n36061), .ALUT(n36062), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2627[11]));
    PFUMX i34306 (.BLUT(n41066), .ALUT(n45209), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2627[4]));
    
endmodule
//
// Verilog Description of module lm32_multiplier
//

module lm32_multiplier (multiplier_result_w, REF_CLK_c, REF_CLK_c_enable_1606, 
            GND_net, VCC_net, operand_1_x, operand_0_x, n45171) /* synthesis syn_module_defined=1 */ ;
    output [31:0]multiplier_result_w;
    input REF_CLK_c;
    input REF_CLK_c_enable_1606;
    input GND_net;
    input VCC_net;
    input [31:0]operand_1_x;
    input [31:0]operand_0_x;
    input n45171;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    wire [63:0]n197;
    
    wire n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, 
        n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, 
        n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, 
        n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, 
        n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, 
        n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, 
        n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, 
        n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, 
        n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, 
        n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, 
        n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, 
        n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, 
        n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, 
        n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, 
        n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, 
        n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, 
        n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, 
        n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, 
        n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, 
        n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, 
        n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, 
        n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, 
        n9019, n9020, n9021, n9022, n9023, n9024, n9025, n8697, 
        n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, 
        n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, 
        n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, 
        n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, 
        n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, 
        n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, 
        n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, 
        n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, 
        n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, 
        n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, 
        n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, 
        n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, 
        n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, 
        n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, 
        n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, 
        n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, 
        n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, 
        n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, 
        n8842;
    
    FD1S3DX result_e3_i0_i0 (.D(n197[0]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[0]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i0.GSR = "ENABLED";
    ALU54B lat_alu_4 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n8879), .SIGNEDIB(n8952), .SIGNEDCIN(n9025), .A35(n8878), 
           .A34(n8877), .A33(n8876), .A32(n8875), .A31(n8874), .A30(n8873), 
           .A29(n8872), .A28(n8871), .A27(n8870), .A26(n8869), .A25(n8868), 
           .A24(n8867), .A23(n8866), .A22(n8865), .A21(n8864), .A20(n8863), 
           .A19(n8862), .A18(n8861), .A17(n8860), .A16(n8859), .A15(n8858), 
           .A14(n8857), .A13(n8856), .A12(n8855), .A11(n8854), .A10(n8853), 
           .A9(n8852), .A8(n8851), .A7(n8850), .A6(n8849), .A5(n8848), 
           .A4(n8847), .A3(n8846), .A2(n8845), .A1(n8844), .A0(n8843), 
           .B35(n8951), .B34(n8950), .B33(n8949), .B32(n8948), .B31(n8947), 
           .B30(n8946), .B29(n8945), .B28(n8944), .B27(n8943), .B26(n8942), 
           .B25(n8941), .B24(n8940), .B23(n8939), .B22(n8938), .B21(n8937), 
           .B20(n8936), .B19(n8935), .B18(n8934), .B17(n8933), .B16(n8932), 
           .B15(n8931), .B14(n8930), .B13(n8929), .B12(n8928), .B11(n8927), 
           .B10(n8926), .B9(n8925), .B8(n8924), .B7(n8923), .B6(n8922), 
           .B5(n8921), .B4(n8920), .B3(n8919), .B2(n8918), .B1(n8917), 
           .B0(n8916), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n8915), .MA34(n8914), .MA33(n8913), .MA32(n8912), .MA31(n8911), 
           .MA30(n8910), .MA29(n8909), .MA28(n8908), .MA27(n8907), .MA26(n8906), 
           .MA25(n8905), .MA24(n8904), .MA23(n8903), .MA22(n8902), .MA21(n8901), 
           .MA20(n8900), .MA19(n8899), .MA18(n8898), .MA17(n8897), .MA16(n8896), 
           .MA15(n8895), .MA14(n8894), .MA13(n8893), .MA12(n8892), .MA11(n8891), 
           .MA10(n8890), .MA9(n8889), .MA8(n8888), .MA7(n8887), .MA6(n8886), 
           .MA5(n8885), .MA4(n8884), .MA3(n8883), .MA2(n8882), .MA1(n8881), 
           .MA0(n8880), .MB35(n8988), .MB34(n8987), .MB33(n8986), .MB32(n8985), 
           .MB31(n8984), .MB30(n8983), .MB29(n8982), .MB28(n8981), .MB27(n8980), 
           .MB26(n8979), .MB25(n8978), .MB24(n8977), .MB23(n8976), .MB22(n8975), 
           .MB21(n8974), .MB20(n8973), .MB19(n8972), .MB18(n8971), .MB17(n8970), 
           .MB16(n8969), .MB15(n8968), .MB14(n8967), .MB13(n8966), .MB12(n8965), 
           .MB11(n8964), .MB10(n8963), .MB9(n8962), .MB8(n8961), .MB7(n8960), 
           .MB6(n8959), .MB5(n8958), .MB4(n8957), .MB3(n8956), .MB2(n8955), 
           .MB1(n8954), .MB0(n8953), .CIN53(n9024), .CIN52(n9023), .CIN51(n9022), 
           .CIN50(n9021), .CIN49(n9020), .CIN48(n9019), .CIN47(n9018), 
           .CIN46(n9017), .CIN45(n9016), .CIN44(n9015), .CIN43(n9014), 
           .CIN42(n9013), .CIN41(n9012), .CIN40(n9011), .CIN39(n9010), 
           .CIN38(n9009), .CIN37(n9008), .CIN36(n9007), .CIN35(n9006), 
           .CIN34(n9005), .CIN33(n9004), .CIN32(n9003), .CIN31(n9002), 
           .CIN30(n9001), .CIN29(n9000), .CIN28(n8999), .CIN27(n8998), 
           .CIN26(n8997), .CIN25(n8996), .CIN24(n8995), .CIN23(n8994), 
           .CIN22(n8993), .CIN21(n8992), .CIN20(n8991), .CIN19(n8990), 
           .CIN18(n8989), .CIN17(n197[17]), .CIN16(n197[16]), .CIN15(n197[15]), 
           .CIN14(n197[14]), .CIN13(n197[13]), .CIN12(n197[12]), .CIN11(n197[11]), 
           .CIN10(n197[10]), .CIN9(n197[9]), .CIN8(n197[8]), .CIN7(n197[7]), 
           .CIN6(n197[6]), .CIN5(n197[5]), .CIN4(n197[4]), .CIN3(n197[3]), 
           .CIN2(n197[2]), .CIN1(n197[1]), .CIN0(n197[0]), .OP10(GND_net), 
           .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), .OP6(GND_net), 
           .OP5(GND_net), .OP4(VCC_net), .OP3(GND_net), .OP2(GND_net), 
           .OP1(GND_net), .OP0(VCC_net), .R13(n197[31]), .R12(n197[30]), 
           .R11(n197[29]), .R10(n197[28]), .R9(n197[27]), .R8(n197[26]), 
           .R7(n197[25]), .R6(n197[24]), .R5(n197[23]), .R4(n197[22]), 
           .R3(n197[21]), .R2(n197[20]), .R1(n197[19]), .R0(n197[18]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam lat_alu_4.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_4.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_4.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_4.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_4.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_4.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_4.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_4.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_4.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_4.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_4.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_4.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_4.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_4.REG_FLAG_CLK = "NONE";
    defparam lat_alu_4.REG_FLAG_CE = "CE0";
    defparam lat_alu_4.REG_FLAG_RST = "RST0";
    defparam lat_alu_4.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_4.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_4.MASK01 = "0x00000000000000";
    defparam lat_alu_4.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_4.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_4.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_4.CLK0_DIV = "ENABLED";
    defparam lat_alu_4.CLK1_DIV = "ENABLED";
    defparam lat_alu_4.CLK2_DIV = "ENABLED";
    defparam lat_alu_4.CLK3_DIV = "ENABLED";
    defparam lat_alu_4.MCPAT = "0x00000000000000";
    defparam lat_alu_4.MASKPAT = "0x00000000000000";
    defparam lat_alu_4.RNDPAT = "0x00000000000000";
    defparam lat_alu_4.GSR = "ENABLED";
    defparam lat_alu_4.RESETMODE = "SYNC";
    defparam lat_alu_4.MULT9_MODE = "DISABLED";
    defparam lat_alu_4.LEGACY = "DISABLED";
    ALU54B lat_alu_3 (.CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
           .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
           .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
           .SIGNEDIA(n8733), .SIGNEDIB(n8806), .SIGNEDCIN(GND_net), .A35(n8732), 
           .A34(n8731), .A33(n8730), .A32(n8729), .A31(n8728), .A30(n8727), 
           .A29(n8726), .A28(n8725), .A27(n8724), .A26(n8723), .A25(n8722), 
           .A24(n8721), .A23(n8720), .A22(n8719), .A21(n8718), .A20(n8717), 
           .A19(n8716), .A18(n8715), .A17(n8714), .A16(n8713), .A15(n8712), 
           .A14(n8711), .A13(n8710), .A12(n8709), .A11(n8708), .A10(n8707), 
           .A9(n8706), .A8(n8705), .A7(n8704), .A6(n8703), .A5(n8702), 
           .A4(n8701), .A3(n8700), .A2(n8699), .A1(n8698), .A0(n8697), 
           .B35(n8805), .B34(n8804), .B33(n8803), .B32(n8802), .B31(n8801), 
           .B30(n8800), .B29(n8799), .B28(n8798), .B27(n8797), .B26(n8796), 
           .B25(n8795), .B24(n8794), .B23(n8793), .B22(n8792), .B21(n8791), 
           .B20(n8790), .B19(n8789), .B18(n8788), .B17(n8787), .B16(n8786), 
           .B15(n8785), .B14(n8784), .B13(n8783), .B12(n8782), .B11(n8781), 
           .B10(n8780), .B9(n8779), .B8(n8778), .B7(n8777), .B6(n8776), 
           .B5(n8775), .B4(n8774), .B3(n8773), .B2(n8772), .B1(n8771), 
           .B0(n8770), .C53(GND_net), .C52(GND_net), .C51(GND_net), 
           .C50(GND_net), .C49(GND_net), .C48(GND_net), .C47(GND_net), 
           .C46(GND_net), .C45(GND_net), .C44(GND_net), .C43(GND_net), 
           .C42(GND_net), .C41(GND_net), .C40(GND_net), .C39(GND_net), 
           .C38(GND_net), .C37(GND_net), .C36(GND_net), .C35(GND_net), 
           .C34(GND_net), .C33(GND_net), .C32(GND_net), .C31(GND_net), 
           .C30(GND_net), .C29(GND_net), .C28(GND_net), .C27(GND_net), 
           .C26(GND_net), .C25(GND_net), .C24(GND_net), .C23(GND_net), 
           .C22(GND_net), .C21(GND_net), .C20(GND_net), .C19(GND_net), 
           .C18(GND_net), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
           .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
           .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
           .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
           .C1(GND_net), .C0(GND_net), .CFB53(GND_net), .CFB52(GND_net), 
           .CFB51(GND_net), .CFB50(GND_net), .CFB49(GND_net), .CFB48(GND_net), 
           .CFB47(GND_net), .CFB46(GND_net), .CFB45(GND_net), .CFB44(GND_net), 
           .CFB43(GND_net), .CFB42(GND_net), .CFB41(GND_net), .CFB40(GND_net), 
           .CFB39(GND_net), .CFB38(GND_net), .CFB37(GND_net), .CFB36(GND_net), 
           .CFB35(GND_net), .CFB34(GND_net), .CFB33(GND_net), .CFB32(GND_net), 
           .CFB31(GND_net), .CFB30(GND_net), .CFB29(GND_net), .CFB28(GND_net), 
           .CFB27(GND_net), .CFB26(GND_net), .CFB25(GND_net), .CFB24(GND_net), 
           .CFB23(GND_net), .CFB22(GND_net), .CFB21(GND_net), .CFB20(GND_net), 
           .CFB19(GND_net), .CFB18(GND_net), .CFB17(GND_net), .CFB16(GND_net), 
           .CFB15(GND_net), .CFB14(GND_net), .CFB13(GND_net), .CFB12(GND_net), 
           .CFB11(GND_net), .CFB10(GND_net), .CFB9(GND_net), .CFB8(GND_net), 
           .CFB7(GND_net), .CFB6(GND_net), .CFB5(GND_net), .CFB4(GND_net), 
           .CFB3(GND_net), .CFB2(GND_net), .CFB1(GND_net), .CFB0(GND_net), 
           .MA35(n8769), .MA34(n8768), .MA33(n8767), .MA32(n8766), .MA31(n8765), 
           .MA30(n8764), .MA29(n8763), .MA28(n8762), .MA27(n8761), .MA26(n8760), 
           .MA25(n8759), .MA24(n8758), .MA23(n8757), .MA22(n8756), .MA21(n8755), 
           .MA20(n8754), .MA19(n8753), .MA18(n8752), .MA17(n8751), .MA16(n8750), 
           .MA15(n8749), .MA14(n8748), .MA13(n8747), .MA12(n8746), .MA11(n8745), 
           .MA10(n8744), .MA9(n8743), .MA8(n8742), .MA7(n8741), .MA6(n8740), 
           .MA5(n8739), .MA4(n8738), .MA3(n8737), .MA2(n8736), .MA1(n8735), 
           .MA0(n8734), .MB35(n8842), .MB34(n8841), .MB33(n8840), .MB32(n8839), 
           .MB31(n8838), .MB30(n8837), .MB29(n8836), .MB28(n8835), .MB27(n8834), 
           .MB26(n8833), .MB25(n8832), .MB24(n8831), .MB23(n8830), .MB22(n8829), 
           .MB21(n8828), .MB20(n8827), .MB19(n8826), .MB18(n8825), .MB17(n8824), 
           .MB16(n8823), .MB15(n8822), .MB14(n8821), .MB13(n8820), .MB12(n8819), 
           .MB11(n8818), .MB10(n8817), .MB9(n8816), .MB8(n8815), .MB7(n8814), 
           .MB6(n8813), .MB5(n8812), .MB4(n8811), .MB3(n8810), .MB2(n8809), 
           .MB1(n8808), .MB0(n8807), .CIN53(GND_net), .CIN52(GND_net), 
           .CIN51(GND_net), .CIN50(GND_net), .CIN49(GND_net), .CIN48(GND_net), 
           .CIN47(GND_net), .CIN46(GND_net), .CIN45(GND_net), .CIN44(GND_net), 
           .CIN43(GND_net), .CIN42(GND_net), .CIN41(GND_net), .CIN40(GND_net), 
           .CIN39(GND_net), .CIN38(GND_net), .CIN37(GND_net), .CIN36(GND_net), 
           .CIN35(GND_net), .CIN34(GND_net), .CIN33(GND_net), .CIN32(GND_net), 
           .CIN31(GND_net), .CIN30(GND_net), .CIN29(GND_net), .CIN28(GND_net), 
           .CIN27(GND_net), .CIN26(GND_net), .CIN25(GND_net), .CIN24(GND_net), 
           .CIN23(GND_net), .CIN22(GND_net), .CIN21(GND_net), .CIN20(GND_net), 
           .CIN19(GND_net), .CIN18(GND_net), .CIN17(GND_net), .CIN16(GND_net), 
           .CIN15(GND_net), .CIN14(GND_net), .CIN13(GND_net), .CIN12(GND_net), 
           .CIN11(GND_net), .CIN10(GND_net), .CIN9(GND_net), .CIN8(GND_net), 
           .CIN7(GND_net), .CIN6(GND_net), .CIN5(GND_net), .CIN4(GND_net), 
           .CIN3(GND_net), .CIN2(GND_net), .CIN1(GND_net), .CIN0(GND_net), 
           .OP10(GND_net), .OP9(VCC_net), .OP8(GND_net), .OP7(GND_net), 
           .OP6(GND_net), .OP5(GND_net), .OP4(GND_net), .OP3(GND_net), 
           .OP2(GND_net), .OP1(GND_net), .OP0(VCC_net), .R53(n9024), 
           .R52(n9023), .R51(n9022), .R50(n9021), .R49(n9020), .R48(n9019), 
           .R47(n9018), .R46(n9017), .R45(n9016), .R44(n9015), .R43(n9014), 
           .R42(n9013), .R41(n9012), .R40(n9011), .R39(n9010), .R38(n9009), 
           .R37(n9008), .R36(n9007), .R35(n9006), .R34(n9005), .R33(n9004), 
           .R32(n9003), .R31(n9002), .R30(n9001), .R29(n9000), .R28(n8999), 
           .R27(n8998), .R26(n8997), .R25(n8996), .R24(n8995), .R23(n8994), 
           .R22(n8993), .R21(n8992), .R20(n8991), .R19(n8990), .R18(n8989), 
           .R17(n197[17]), .R16(n197[16]), .R15(n197[15]), .R14(n197[14]), 
           .R13(n197[13]), .R12(n197[12]), .R11(n197[11]), .R10(n197[10]), 
           .R9(n197[9]), .R8(n197[8]), .R7(n197[7]), .R6(n197[6]), .R5(n197[5]), 
           .R4(n197[4]), .R3(n197[3]), .R2(n197[2]), .R1(n197[1]), .R0(n197[0]), 
           .SIGNEDR(n9025));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam lat_alu_3.REG_INPUTC0_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTC0_CE = "CE0";
    defparam lat_alu_3.REG_INPUTC0_RST = "RST0";
    defparam lat_alu_3.REG_INPUTC1_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTC1_CE = "CE0";
    defparam lat_alu_3.REG_INPUTC1_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP0_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_0_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEOP0_0_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP1_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEOP0_1_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEOP0_1_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEOP1_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_0_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_0_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEIN_0_RST = "RST0";
    defparam lat_alu_3.REG_OPCODEIN_1_CLK = "NONE";
    defparam lat_alu_3.REG_OPCODEIN_1_CE = "CE0";
    defparam lat_alu_3.REG_OPCODEIN_1_RST = "RST0";
    defparam lat_alu_3.REG_OUTPUT0_CLK = "NONE";
    defparam lat_alu_3.REG_OUTPUT0_CE = "CE0";
    defparam lat_alu_3.REG_OUTPUT0_RST = "RST0";
    defparam lat_alu_3.REG_OUTPUT1_CLK = "NONE";
    defparam lat_alu_3.REG_OUTPUT1_CE = "CE0";
    defparam lat_alu_3.REG_OUTPUT1_RST = "RST0";
    defparam lat_alu_3.REG_FLAG_CLK = "NONE";
    defparam lat_alu_3.REG_FLAG_CE = "CE0";
    defparam lat_alu_3.REG_FLAG_RST = "RST0";
    defparam lat_alu_3.MCPAT_SOURCE = "STATIC";
    defparam lat_alu_3.MASKPAT_SOURCE = "STATIC";
    defparam lat_alu_3.MASK01 = "0x00000000000000";
    defparam lat_alu_3.REG_INPUTCFB_CLK = "NONE";
    defparam lat_alu_3.REG_INPUTCFB_CE = "CE0";
    defparam lat_alu_3.REG_INPUTCFB_RST = "RST0";
    defparam lat_alu_3.CLK0_DIV = "ENABLED";
    defparam lat_alu_3.CLK1_DIV = "ENABLED";
    defparam lat_alu_3.CLK2_DIV = "ENABLED";
    defparam lat_alu_3.CLK3_DIV = "ENABLED";
    defparam lat_alu_3.MCPAT = "0x00000000000000";
    defparam lat_alu_3.MASKPAT = "0x00000000000000";
    defparam lat_alu_3.RNDPAT = "0x00000000000000";
    defparam lat_alu_3.GSR = "ENABLED";
    defparam lat_alu_3.RESETMODE = "SYNC";
    defparam lat_alu_3.MULT9_MODE = "DISABLED";
    defparam lat_alu_3.LEGACY = "DISABLED";
    MULT18X18D lat_mult_2 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(operand_1_x[31]), .A12(operand_1_x[30]), 
            .A11(operand_1_x[29]), .A10(operand_1_x[28]), .A9(operand_1_x[27]), 
            .A8(operand_1_x[26]), .A7(operand_1_x[25]), .A6(operand_1_x[24]), 
            .A5(operand_1_x[23]), .A4(operand_1_x[22]), .A3(operand_1_x[21]), 
            .A2(operand_1_x[20]), .A1(operand_1_x[19]), .A0(operand_1_x[18]), 
            .B17(GND_net), .B16(GND_net), .B15(GND_net), .B14(GND_net), 
            .B13(operand_0_x[31]), .B12(operand_0_x[30]), .B11(operand_0_x[29]), 
            .B10(operand_0_x[28]), .B9(operand_0_x[27]), .B8(operand_0_x[26]), 
            .B7(operand_0_x[25]), .B6(operand_0_x[24]), .B5(operand_0_x[23]), 
            .B4(operand_0_x[22]), .B3(operand_0_x[21]), .B2(operand_0_x[20]), 
            .B1(operand_0_x[19]), .B0(operand_0_x[18]), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(REF_CLK_c), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(n45171), .CE2(GND_net), .CE1(GND_net), 
            .CE0(VCC_net), .RST3(REF_CLK_c_enable_1606), .RST2(GND_net), 
            .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), 
            .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), 
            .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), 
            .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), 
            .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), 
            .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), 
            .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), 
            .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), 
            .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), 
            .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n8933), .ROA16(n8932), 
            .ROA15(n8931), .ROA14(n8930), .ROA13(n8929), .ROA12(n8928), 
            .ROA11(n8927), .ROA10(n8926), .ROA9(n8925), .ROA8(n8924), 
            .ROA7(n8923), .ROA6(n8922), .ROA5(n8921), .ROA4(n8920), 
            .ROA3(n8919), .ROA2(n8918), .ROA1(n8917), .ROA0(n8916), 
            .ROB17(n8951), .ROB16(n8950), .ROB15(n8949), .ROB14(n8948), 
            .ROB13(n8947), .ROB12(n8946), .ROB11(n8945), .ROB10(n8944), 
            .ROB9(n8943), .ROB8(n8942), .ROB7(n8941), .ROB6(n8940), 
            .ROB5(n8939), .ROB4(n8938), .ROB3(n8937), .ROB2(n8936), 
            .ROB1(n8935), .ROB0(n8934), .P35(n8988), .P34(n8987), .P33(n8986), 
            .P32(n8985), .P31(n8984), .P30(n8983), .P29(n8982), .P28(n8981), 
            .P27(n8980), .P26(n8979), .P25(n8978), .P24(n8977), .P23(n8976), 
            .P22(n8975), .P21(n8974), .P20(n8973), .P19(n8972), .P18(n8971), 
            .P17(n8970), .P16(n8969), .P15(n8968), .P14(n8967), .P13(n8966), 
            .P12(n8965), .P11(n8964), .P10(n8963), .P9(n8962), .P8(n8961), 
            .P7(n8960), .P6(n8959), .P5(n8958), .P4(n8957), .P3(n8956), 
            .P2(n8955), .P1(n8954), .P0(n8953), .SIGNEDP(n8952));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam lat_mult_2.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_2.REG_INPUTA_CE = "CE3";
    defparam lat_mult_2.REG_INPUTA_RST = "RST3";
    defparam lat_mult_2.REG_INPUTB_CLK = "CLK3";
    defparam lat_mult_2.REG_INPUTB_CE = "CE3";
    defparam lat_mult_2.REG_INPUTB_RST = "RST3";
    defparam lat_mult_2.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_2.REG_INPUTC_CE = "CE0";
    defparam lat_mult_2.REG_INPUTC_RST = "RST0";
    defparam lat_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_2.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_2.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_2.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_2.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_2.CLK0_DIV = "ENABLED";
    defparam lat_mult_2.CLK1_DIV = "ENABLED";
    defparam lat_mult_2.CLK2_DIV = "ENABLED";
    defparam lat_mult_2.CLK3_DIV = "ENABLED";
    defparam lat_mult_2.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_2.GSR = "ENABLED";
    defparam lat_mult_2.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_2.MULT_BYPASS = "DISABLED";
    defparam lat_mult_2.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_1 (.A17(operand_1_x[17]), .A16(operand_1_x[16]), 
            .A15(operand_1_x[15]), .A14(operand_1_x[14]), .A13(operand_1_x[13]), 
            .A12(operand_1_x[12]), .A11(operand_1_x[11]), .A10(operand_1_x[10]), 
            .A9(operand_1_x[9]), .A8(operand_1_x[8]), .A7(operand_1_x[7]), 
            .A6(operand_1_x[6]), .A5(operand_1_x[5]), .A4(operand_1_x[4]), 
            .A3(operand_1_x[3]), .A2(operand_1_x[2]), .A1(operand_1_x[1]), 
            .A0(operand_1_x[0]), .B17(GND_net), .B16(GND_net), .B15(GND_net), 
            .B14(GND_net), .B13(operand_0_x[31]), .B12(operand_0_x[30]), 
            .B11(operand_0_x[29]), .B10(operand_0_x[28]), .B9(operand_0_x[27]), 
            .B8(operand_0_x[26]), .B7(operand_0_x[25]), .B6(operand_0_x[24]), 
            .B5(operand_0_x[23]), .B4(operand_0_x[22]), .B3(operand_0_x[21]), 
            .B2(operand_0_x[20]), .B1(operand_0_x[19]), .B0(operand_0_x[18]), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(REF_CLK_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(n45171), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(REF_CLK_c_enable_1606), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n8860), 
            .ROA16(n8859), .ROA15(n8858), .ROA14(n8857), .ROA13(n8856), 
            .ROA12(n8855), .ROA11(n8854), .ROA10(n8853), .ROA9(n8852), 
            .ROA8(n8851), .ROA7(n8850), .ROA6(n8849), .ROA5(n8848), 
            .ROA4(n8847), .ROA3(n8846), .ROA2(n8845), .ROA1(n8844), 
            .ROA0(n8843), .ROB17(n8878), .ROB16(n8877), .ROB15(n8876), 
            .ROB14(n8875), .ROB13(n8874), .ROB12(n8873), .ROB11(n8872), 
            .ROB10(n8871), .ROB9(n8870), .ROB8(n8869), .ROB7(n8868), 
            .ROB6(n8867), .ROB5(n8866), .ROB4(n8865), .ROB3(n8864), 
            .ROB2(n8863), .ROB1(n8862), .ROB0(n8861), .P35(n8915), .P34(n8914), 
            .P33(n8913), .P32(n8912), .P31(n8911), .P30(n8910), .P29(n8909), 
            .P28(n8908), .P27(n8907), .P26(n8906), .P25(n8905), .P24(n8904), 
            .P23(n8903), .P22(n8902), .P21(n8901), .P20(n8900), .P19(n8899), 
            .P18(n8898), .P17(n8897), .P16(n8896), .P15(n8895), .P14(n8894), 
            .P13(n8893), .P12(n8892), .P11(n8891), .P10(n8890), .P9(n8889), 
            .P8(n8888), .P7(n8887), .P6(n8886), .P5(n8885), .P4(n8884), 
            .P3(n8883), .P2(n8882), .P1(n8881), .P0(n8880), .SIGNEDP(n8879));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam lat_mult_1.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_1.REG_INPUTA_CE = "CE3";
    defparam lat_mult_1.REG_INPUTA_RST = "RST3";
    defparam lat_mult_1.REG_INPUTB_CLK = "CLK3";
    defparam lat_mult_1.REG_INPUTB_CE = "CE3";
    defparam lat_mult_1.REG_INPUTB_RST = "RST3";
    defparam lat_mult_1.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_1.REG_INPUTC_CE = "CE0";
    defparam lat_mult_1.REG_INPUTC_RST = "RST0";
    defparam lat_mult_1.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_1.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_1.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_1.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_1.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_1.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_1.CLK0_DIV = "ENABLED";
    defparam lat_mult_1.CLK1_DIV = "ENABLED";
    defparam lat_mult_1.CLK2_DIV = "ENABLED";
    defparam lat_mult_1.CLK3_DIV = "ENABLED";
    defparam lat_mult_1.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_1.GSR = "ENABLED";
    defparam lat_mult_1.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_1.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_1.MULT_BYPASS = "DISABLED";
    defparam lat_mult_1.RESETMODE = "ASYNC";
    MULT18X18D lat_mult_0 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(operand_1_x[31]), .A12(operand_1_x[30]), 
            .A11(operand_1_x[29]), .A10(operand_1_x[28]), .A9(operand_1_x[27]), 
            .A8(operand_1_x[26]), .A7(operand_1_x[25]), .A6(operand_1_x[24]), 
            .A5(operand_1_x[23]), .A4(operand_1_x[22]), .A3(operand_1_x[21]), 
            .A2(operand_1_x[20]), .A1(operand_1_x[19]), .A0(operand_1_x[18]), 
            .B17(operand_0_x[17]), .B16(operand_0_x[16]), .B15(operand_0_x[15]), 
            .B14(operand_0_x[14]), .B13(operand_0_x[13]), .B12(operand_0_x[12]), 
            .B11(operand_0_x[11]), .B10(operand_0_x[10]), .B9(operand_0_x[9]), 
            .B8(operand_0_x[8]), .B7(operand_0_x[7]), .B6(operand_0_x[6]), 
            .B5(operand_0_x[5]), .B4(operand_0_x[4]), .B3(operand_0_x[3]), 
            .B2(operand_0_x[2]), .B1(operand_0_x[1]), .B0(operand_0_x[0]), 
            .C17(GND_net), .C16(GND_net), .C15(GND_net), .C14(GND_net), 
            .C13(GND_net), .C12(GND_net), .C11(GND_net), .C10(GND_net), 
            .C9(GND_net), .C8(GND_net), .C7(GND_net), .C6(GND_net), 
            .C5(GND_net), .C4(GND_net), .C3(GND_net), .C2(GND_net), 
            .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), .SIGNEDB(GND_net), 
            .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(REF_CLK_c), .CLK2(GND_net), 
            .CLK1(GND_net), .CLK0(GND_net), .CE3(n45171), .CE2(GND_net), 
            .CE1(GND_net), .CE0(VCC_net), .RST3(REF_CLK_c_enable_1606), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n8787), 
            .ROA16(n8786), .ROA15(n8785), .ROA14(n8784), .ROA13(n8783), 
            .ROA12(n8782), .ROA11(n8781), .ROA10(n8780), .ROA9(n8779), 
            .ROA8(n8778), .ROA7(n8777), .ROA6(n8776), .ROA5(n8775), 
            .ROA4(n8774), .ROA3(n8773), .ROA2(n8772), .ROA1(n8771), 
            .ROA0(n8770), .ROB17(n8805), .ROB16(n8804), .ROB15(n8803), 
            .ROB14(n8802), .ROB13(n8801), .ROB12(n8800), .ROB11(n8799), 
            .ROB10(n8798), .ROB9(n8797), .ROB8(n8796), .ROB7(n8795), 
            .ROB6(n8794), .ROB5(n8793), .ROB4(n8792), .ROB3(n8791), 
            .ROB2(n8790), .ROB1(n8789), .ROB0(n8788), .P35(n8842), .P34(n8841), 
            .P33(n8840), .P32(n8839), .P31(n8838), .P30(n8837), .P29(n8836), 
            .P28(n8835), .P27(n8834), .P26(n8833), .P25(n8832), .P24(n8831), 
            .P23(n8830), .P22(n8829), .P21(n8828), .P20(n8827), .P19(n8826), 
            .P18(n8825), .P17(n8824), .P16(n8823), .P15(n8822), .P14(n8821), 
            .P13(n8820), .P12(n8819), .P11(n8818), .P10(n8817), .P9(n8816), 
            .P8(n8815), .P7(n8814), .P6(n8813), .P5(n8812), .P4(n8811), 
            .P3(n8810), .P2(n8809), .P1(n8808), .P0(n8807), .SIGNEDP(n8806));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam lat_mult_0.REG_INPUTA_CLK = "CLK3";
    defparam lat_mult_0.REG_INPUTA_CE = "CE3";
    defparam lat_mult_0.REG_INPUTA_RST = "RST3";
    defparam lat_mult_0.REG_INPUTB_CLK = "CLK3";
    defparam lat_mult_0.REG_INPUTB_CE = "CE3";
    defparam lat_mult_0.REG_INPUTB_RST = "RST3";
    defparam lat_mult_0.REG_INPUTC_CLK = "NONE";
    defparam lat_mult_0.REG_INPUTC_CE = "CE0";
    defparam lat_mult_0.REG_INPUTC_RST = "RST0";
    defparam lat_mult_0.REG_PIPELINE_CLK = "NONE";
    defparam lat_mult_0.REG_PIPELINE_CE = "CE0";
    defparam lat_mult_0.REG_PIPELINE_RST = "RST0";
    defparam lat_mult_0.REG_OUTPUT_CLK = "NONE";
    defparam lat_mult_0.REG_OUTPUT_CE = "CE0";
    defparam lat_mult_0.REG_OUTPUT_RST = "RST0";
    defparam lat_mult_0.CLK0_DIV = "ENABLED";
    defparam lat_mult_0.CLK1_DIV = "ENABLED";
    defparam lat_mult_0.CLK2_DIV = "ENABLED";
    defparam lat_mult_0.CLK3_DIV = "ENABLED";
    defparam lat_mult_0.HIGHSPEED_CLK = "NONE";
    defparam lat_mult_0.GSR = "ENABLED";
    defparam lat_mult_0.CAS_MATCH_REG = "FALSE";
    defparam lat_mult_0.SOURCEB_MODE = "B_SHIFT";
    defparam lat_mult_0.MULT_BYPASS = "DISABLED";
    defparam lat_mult_0.RESETMODE = "ASYNC";
    MULT18X18D result_mult_2 (.A17(operand_1_x[17]), .A16(operand_1_x[16]), 
            .A15(operand_1_x[15]), .A14(operand_1_x[14]), .A13(operand_1_x[13]), 
            .A12(operand_1_x[12]), .A11(operand_1_x[11]), .A10(operand_1_x[10]), 
            .A9(operand_1_x[9]), .A8(operand_1_x[8]), .A7(operand_1_x[7]), 
            .A6(operand_1_x[6]), .A5(operand_1_x[5]), .A4(operand_1_x[4]), 
            .A3(operand_1_x[3]), .A2(operand_1_x[2]), .A1(operand_1_x[1]), 
            .A0(operand_1_x[0]), .B17(operand_0_x[17]), .B16(operand_0_x[16]), 
            .B15(operand_0_x[15]), .B14(operand_0_x[14]), .B13(operand_0_x[13]), 
            .B12(operand_0_x[12]), .B11(operand_0_x[11]), .B10(operand_0_x[10]), 
            .B9(operand_0_x[9]), .B8(operand_0_x[8]), .B7(operand_0_x[7]), 
            .B6(operand_0_x[6]), .B5(operand_0_x[5]), .B4(operand_0_x[4]), 
            .B3(operand_0_x[3]), .B2(operand_0_x[2]), .B1(operand_0_x[1]), 
            .B0(operand_0_x[0]), .C17(GND_net), .C16(GND_net), .C15(GND_net), 
            .C14(GND_net), .C13(GND_net), .C12(GND_net), .C11(GND_net), 
            .C10(GND_net), .C9(GND_net), .C8(GND_net), .C7(GND_net), 
            .C6(GND_net), .C5(GND_net), .C4(GND_net), .C3(GND_net), 
            .C2(GND_net), .C1(GND_net), .C0(GND_net), .SIGNEDA(GND_net), 
            .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), .CLK3(REF_CLK_c), 
            .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), .CE3(n45171), 
            .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), .RST3(REF_CLK_c_enable_1606), 
            .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), .SRIA17(GND_net), 
            .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), .SRIA13(GND_net), 
            .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), .SRIA9(GND_net), 
            .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), .SRIA5(GND_net), 
            .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), .SRIA1(GND_net), 
            .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), .SRIB15(GND_net), 
            .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), .SRIB11(GND_net), 
            .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), .SRIB7(GND_net), 
            .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), .SRIB3(GND_net), 
            .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), .ROA17(n8714), 
            .ROA16(n8713), .ROA15(n8712), .ROA14(n8711), .ROA13(n8710), 
            .ROA12(n8709), .ROA11(n8708), .ROA10(n8707), .ROA9(n8706), 
            .ROA8(n8705), .ROA7(n8704), .ROA6(n8703), .ROA5(n8702), 
            .ROA4(n8701), .ROA3(n8700), .ROA2(n8699), .ROA1(n8698), 
            .ROA0(n8697), .ROB17(n8732), .ROB16(n8731), .ROB15(n8730), 
            .ROB14(n8729), .ROB13(n8728), .ROB12(n8727), .ROB11(n8726), 
            .ROB10(n8725), .ROB9(n8724), .ROB8(n8723), .ROB7(n8722), 
            .ROB6(n8721), .ROB5(n8720), .ROB4(n8719), .ROB3(n8718), 
            .ROB2(n8717), .ROB1(n8716), .ROB0(n8715), .P35(n8769), .P34(n8768), 
            .P33(n8767), .P32(n8766), .P31(n8765), .P30(n8764), .P29(n8763), 
            .P28(n8762), .P27(n8761), .P26(n8760), .P25(n8759), .P24(n8758), 
            .P23(n8757), .P22(n8756), .P21(n8755), .P20(n8754), .P19(n8753), 
            .P18(n8752), .P17(n8751), .P16(n8750), .P15(n8749), .P14(n8748), 
            .P13(n8747), .P12(n8746), .P11(n8745), .P10(n8744), .P9(n8743), 
            .P8(n8742), .P7(n8741), .P6(n8740), .P5(n8739), .P4(n8738), 
            .P3(n8737), .P2(n8736), .P1(n8735), .P0(n8734), .SIGNEDP(n8733));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_mult_2.REG_INPUTA_CLK = "CLK3";
    defparam result_mult_2.REG_INPUTA_CE = "CE3";
    defparam result_mult_2.REG_INPUTA_RST = "RST3";
    defparam result_mult_2.REG_INPUTB_CLK = "CLK3";
    defparam result_mult_2.REG_INPUTB_CE = "CE3";
    defparam result_mult_2.REG_INPUTB_RST = "RST3";
    defparam result_mult_2.REG_INPUTC_CLK = "NONE";
    defparam result_mult_2.REG_INPUTC_CE = "CE0";
    defparam result_mult_2.REG_INPUTC_RST = "RST0";
    defparam result_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam result_mult_2.REG_PIPELINE_CE = "CE0";
    defparam result_mult_2.REG_PIPELINE_RST = "RST0";
    defparam result_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam result_mult_2.REG_OUTPUT_CE = "CE0";
    defparam result_mult_2.REG_OUTPUT_RST = "RST0";
    defparam result_mult_2.CLK0_DIV = "ENABLED";
    defparam result_mult_2.CLK1_DIV = "ENABLED";
    defparam result_mult_2.CLK2_DIV = "ENABLED";
    defparam result_mult_2.CLK3_DIV = "ENABLED";
    defparam result_mult_2.HIGHSPEED_CLK = "NONE";
    defparam result_mult_2.GSR = "ENABLED";
    defparam result_mult_2.CAS_MATCH_REG = "FALSE";
    defparam result_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam result_mult_2.MULT_BYPASS = "DISABLED";
    defparam result_mult_2.RESETMODE = "ASYNC";
    FD1S3DX result_e3_i0_i1 (.D(n197[1]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[1]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i1.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i2 (.D(n197[2]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[2]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i2.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i3 (.D(n197[3]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[3]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i3.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i4 (.D(n197[4]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[4]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i4.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i5 (.D(n197[5]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[5]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i5.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i6 (.D(n197[6]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[6]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i6.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i7 (.D(n197[7]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[7]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i7.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i8 (.D(n197[8]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[8]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i8.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i9 (.D(n197[9]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[9]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i9.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i10 (.D(n197[10]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[10]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i10.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i11 (.D(n197[11]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[11]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i11.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i12 (.D(n197[12]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[12]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i12.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i13 (.D(n197[13]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[13]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i13.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i14 (.D(n197[14]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[14]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i14.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i15 (.D(n197[15]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[15]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i15.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i16 (.D(n197[16]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[16]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i16.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i17 (.D(n197[17]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[17]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i17.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i18 (.D(n197[18]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[18]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i18.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i19 (.D(n197[19]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[19]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i19.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i20 (.D(n197[20]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[20]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i20.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i21 (.D(n197[21]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[21]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i21.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i22 (.D(n197[22]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[22]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i22.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i23 (.D(n197[23]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[23]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i23.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i24 (.D(n197[24]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[24]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i24.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i25 (.D(n197[25]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[25]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i25.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i26 (.D(n197[26]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[26]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i26.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i27 (.D(n197[27]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[27]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i27.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i28 (.D(n197[28]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[28]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i28.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i29 (.D(n197[29]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[29]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i29.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i30 (.D(n197[30]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[30]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i30.GSR = "ENABLED";
    FD1S3DX result_e3_i0_i31 (.D(n197[31]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(multiplier_result_w[31]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    defparam result_e3_i0_i31.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module lm32_mc_arithmetic
//

module lm32_mc_arithmetic (REF_CLK_c, REF_CLK_c_enable_1606, b, REF_CLK_c_enable_1366, 
            d_result_1, p, mc_result_x, divide_by_zero_x, cycles_5__N_2934, 
            \a[31] , GND_net, VCC_net, n32636, n15, n41231, n45183, 
            t, d_result_0, n45181, n41216, n41196, q_d, n32608, 
            n41197, n20863, n32652) /* synthesis syn_module_defined=1 */ ;
    input REF_CLK_c;
    input REF_CLK_c_enable_1606;
    output [31:0]b;
    input REF_CLK_c_enable_1366;
    input [31:0]d_result_1;
    output [31:0]p;
    output [31:0]mc_result_x;
    output divide_by_zero_x;
    output cycles_5__N_2934;
    output \a[31] ;
    input GND_net;
    input VCC_net;
    input n32636;
    input n15;
    input n41231;
    input n45183;
    input [32:0]t;
    input [31:0]d_result_0;
    input n45181;
    input n41216;
    input n41196;
    input q_d;
    input n32608;
    input n41197;
    input n20863;
    input n32652;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    
    wire cycles_5__N_2936, n9349;
    wire [31:0]p_31__N_2829;
    wire [31:0]a;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(133[22:23])
    wire [31:0]a_31__N_2861;
    wire [31:0]result_x_31__N_2797;
    
    wire divide_by_zero_x_N_3086;
    wire [5:0]cycles;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(140[11:17])
    wire [5:0]cycles_5__N_2928;
    
    wire n41445, n41396, n1;
    wire [2:0]state;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(139[26:31])
    
    wire n9351, n9353;
    wire [31:0]p_c;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(132[22:23])
    
    wire n35552, n31889, n31888, n31887, n31886, n35551, n31881, 
        n31880, n31879, n31878, n31885, n31884, n31883, n31882, 
        n35550, n31873, n31872, n31871, n31870, n31877, n31876, 
        n31875, n31874, n35549, n31865, n31864, n31863, n31862, 
        n31869, n31868, n31867, n31866, n31858, n31861, n31860, 
        n31859, divide_by_zero_x_N_3090, n35380, n9312, n1_adj_6104, 
        n1_adj_6105, n1_adj_6106, n1_adj_6107, n1_adj_6108, n1_adj_6109, 
        n1_adj_6110, n1_adj_6111, n1_adj_6112, n1_adj_6113, n1_adj_6114, 
        n1_adj_6115, n1_adj_6116, n1_adj_6117, n1_adj_6118, n1_adj_6119, 
        n1_adj_6120, n1_adj_6121, n1_adj_6122, n1_adj_6123, n1_adj_6124, 
        n1_adj_6125, n1_adj_6126, n1_adj_6127, n1_adj_6128, n1_adj_6129, 
        n1_adj_6130, n1_adj_6131, n1_adj_6132, n1_adj_6133, n1_adj_6134, 
        n1_adj_6135, n1_adj_6136;
    wire [31:0]a_31__N_3014;
    
    wire n1_adj_6137, n1_adj_6138, n2, n4, n1_adj_6139, n2_adj_6140, 
        n1_adj_6141, n2_adj_6142, n1_adj_6143, n2_adj_6144, n1_adj_6145, 
        n2_adj_6146, n1_adj_6147, n2_adj_6148, n1_adj_6149, n2_adj_6150, 
        n1_adj_6151, n2_adj_6152, n1_adj_6153, n2_adj_6154, n1_adj_6155, 
        n2_adj_6156, n4_adj_6157, n1_adj_6158, n2_adj_6159, n4_adj_6160, 
        n1_adj_6161, n2_adj_6162, n1_adj_6163, n2_adj_6164, n4_adj_6165, 
        n1_adj_6166, n2_adj_6167, n1_adj_6168, n2_adj_6169, n4_adj_6170, 
        n1_adj_6171, n2_adj_6172, n1_adj_6173, n2_adj_6174, n1_adj_6175, 
        n2_adj_6176, n4_adj_6177, n1_adj_6178, n2_adj_6179, n1_adj_6180, 
        n2_adj_6181, n1_adj_6182, n2_adj_6183, n4_adj_6184, n4_adj_6185, 
        n4_adj_6186, n1_adj_6187, n2_adj_6188, n1_adj_6189, n2_adj_6190, 
        n1_adj_6191, n1_adj_6192, n41293, n41378, n32614, n32658;
    
    FD1S3DX state_FSM_i1 (.D(n9349), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(cycles_5__N_2936));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam state_FSM_i1.GSR = "ENABLED";
    FD1P3DX b_i0_i0 (.D(d_result_1[0]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i0.GSR = "ENABLED";
    FD1S3DX p_i0 (.D(p_31__N_2829[0]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i0.GSR = "ENABLED";
    FD1S3DX a_i0 (.D(a_31__N_2861[0]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0.GSR = "ENABLED";
    FD1S3DX result_x_i0 (.D(result_x_31__N_2797[0]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0.GSR = "ENABLED";
    FD1S3DX divide_by_zero_x_58 (.D(divide_by_zero_x_N_3086), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(divide_by_zero_x)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam divide_by_zero_x_58.GSR = "ENABLED";
    FD1S3DX cycles_i0 (.D(cycles_5__N_2928[0]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(cycles[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam cycles_i0.GSR = "ENABLED";
    LUT4 select_1205_Select_3_i1_3_lut_4_lut (.A(cycles[2]), .B(n41445), 
         .C(n41396), .D(cycles[3]), .Z(n1)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B !((D)+!C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(250[26:39])
    defparam select_1205_Select_3_i1_3_lut_4_lut.init = 16'he010;
    FD1S3DX state_FSM_i2 (.D(n9351), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(state[0]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam state_FSM_i2.GSR = "ENABLED";
    FD1S3BX state_FSM_i3 (.D(n9353), .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), 
            .Q(cycles_5__N_2934));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam state_FSM_i3.GSR = "ENABLED";
    FD1P3DX b_i0_i1 (.D(d_result_1[1]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i1.GSR = "ENABLED";
    FD1P3DX b_i0_i2 (.D(d_result_1[2]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i2.GSR = "ENABLED";
    FD1P3DX b_i0_i3 (.D(d_result_1[3]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i3.GSR = "ENABLED";
    FD1P3DX b_i0_i4 (.D(d_result_1[4]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i4.GSR = "ENABLED";
    FD1P3DX b_i0_i5 (.D(d_result_1[5]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i5.GSR = "ENABLED";
    FD1P3DX b_i0_i6 (.D(d_result_1[6]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i6.GSR = "ENABLED";
    FD1P3DX b_i0_i7 (.D(d_result_1[7]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i7.GSR = "ENABLED";
    FD1P3DX b_i0_i8 (.D(d_result_1[8]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i8.GSR = "ENABLED";
    FD1P3DX b_i0_i9 (.D(d_result_1[9]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i9.GSR = "ENABLED";
    FD1P3DX b_i0_i10 (.D(d_result_1[10]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i10.GSR = "ENABLED";
    FD1P3DX b_i0_i11 (.D(d_result_1[11]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i11.GSR = "ENABLED";
    FD1P3DX b_i0_i12 (.D(d_result_1[12]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i12.GSR = "ENABLED";
    FD1P3DX b_i0_i13 (.D(d_result_1[13]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i13.GSR = "ENABLED";
    FD1P3DX b_i0_i14 (.D(d_result_1[14]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i14.GSR = "ENABLED";
    FD1P3DX b_i0_i15 (.D(d_result_1[15]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i15.GSR = "ENABLED";
    FD1P3DX b_i0_i16 (.D(d_result_1[16]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i16.GSR = "ENABLED";
    FD1P3DX b_i0_i17 (.D(d_result_1[17]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i17.GSR = "ENABLED";
    FD1P3DX b_i0_i18 (.D(d_result_1[18]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i18.GSR = "ENABLED";
    FD1P3DX b_i0_i19 (.D(d_result_1[19]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i19.GSR = "ENABLED";
    FD1P3DX b_i0_i20 (.D(d_result_1[20]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i20.GSR = "ENABLED";
    FD1P3DX b_i0_i21 (.D(d_result_1[21]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i21.GSR = "ENABLED";
    FD1P3DX b_i0_i22 (.D(d_result_1[22]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i22.GSR = "ENABLED";
    FD1P3DX b_i0_i23 (.D(d_result_1[23]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i23.GSR = "ENABLED";
    FD1P3DX b_i0_i24 (.D(d_result_1[24]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i24.GSR = "ENABLED";
    FD1P3DX b_i0_i25 (.D(d_result_1[25]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i25.GSR = "ENABLED";
    FD1P3DX b_i0_i26 (.D(d_result_1[26]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i26.GSR = "ENABLED";
    FD1P3DX b_i0_i27 (.D(d_result_1[27]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i27.GSR = "ENABLED";
    FD1P3DX b_i0_i28 (.D(d_result_1[28]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i28.GSR = "ENABLED";
    FD1P3DX b_i0_i29 (.D(d_result_1[29]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i29.GSR = "ENABLED";
    FD1P3DX b_i0_i30 (.D(d_result_1[30]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i30.GSR = "ENABLED";
    FD1P3DX b_i0_i31 (.D(d_result_1[31]), .SP(REF_CLK_c_enable_1366), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(b[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b_i0_i31.GSR = "ENABLED";
    FD1S3DX p_i1 (.D(p_31__N_2829[1]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i1.GSR = "ENABLED";
    FD1S3DX p_i2 (.D(p_31__N_2829[2]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i2.GSR = "ENABLED";
    FD1S3DX p_i3 (.D(p_31__N_2829[3]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i3.GSR = "ENABLED";
    FD1S3DX p_i4 (.D(p_31__N_2829[4]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i4.GSR = "ENABLED";
    FD1S3DX p_i5 (.D(p_31__N_2829[5]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i5.GSR = "ENABLED";
    FD1S3DX p_i6 (.D(p_31__N_2829[6]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i6.GSR = "ENABLED";
    FD1S3DX p_i7 (.D(p_31__N_2829[7]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i7.GSR = "ENABLED";
    FD1S3DX p_i8 (.D(p_31__N_2829[8]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i8.GSR = "ENABLED";
    FD1S3DX p_i9 (.D(p_31__N_2829[9]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i9.GSR = "ENABLED";
    FD1S3DX p_i10 (.D(p_31__N_2829[10]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i10.GSR = "ENABLED";
    FD1S3DX p_i11 (.D(p_31__N_2829[11]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i11.GSR = "ENABLED";
    FD1S3DX p_i12 (.D(p_31__N_2829[12]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i12.GSR = "ENABLED";
    FD1S3DX p_i13 (.D(p_31__N_2829[13]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i13.GSR = "ENABLED";
    FD1S3DX p_i14 (.D(p_31__N_2829[14]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i14.GSR = "ENABLED";
    FD1S3DX p_i15 (.D(p_31__N_2829[15]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i15.GSR = "ENABLED";
    FD1S3DX p_i16 (.D(p_31__N_2829[16]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i16.GSR = "ENABLED";
    FD1S3DX p_i17 (.D(p_31__N_2829[17]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i17.GSR = "ENABLED";
    FD1S3DX p_i18 (.D(p_31__N_2829[18]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i18.GSR = "ENABLED";
    FD1S3DX p_i19 (.D(p_31__N_2829[19]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i19.GSR = "ENABLED";
    FD1S3DX p_i20 (.D(p_31__N_2829[20]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i20.GSR = "ENABLED";
    FD1S3DX p_i21 (.D(p_31__N_2829[21]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i21.GSR = "ENABLED";
    FD1S3DX p_i22 (.D(p_31__N_2829[22]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i22.GSR = "ENABLED";
    FD1S3DX p_i23 (.D(p_31__N_2829[23]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i23.GSR = "ENABLED";
    FD1S3DX p_i24 (.D(p_31__N_2829[24]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i24.GSR = "ENABLED";
    FD1S3DX p_i25 (.D(p_31__N_2829[25]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i25.GSR = "ENABLED";
    FD1S3DX p_i26 (.D(p_31__N_2829[26]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i26.GSR = "ENABLED";
    FD1S3DX p_i27 (.D(p_31__N_2829[27]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i27.GSR = "ENABLED";
    FD1S3DX p_i28 (.D(p_31__N_2829[28]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i28.GSR = "ENABLED";
    FD1S3DX p_i29 (.D(p_31__N_2829[29]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i29.GSR = "ENABLED";
    FD1S3DX p_i30 (.D(p_31__N_2829[30]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i30.GSR = "ENABLED";
    FD1S3DX p_i31 (.D(p_31__N_2829[31]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(p_c[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p_i31.GSR = "ENABLED";
    FD1S3DX a_i1 (.D(a_31__N_2861[1]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i1.GSR = "ENABLED";
    FD1S3DX a_i2 (.D(a_31__N_2861[2]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i2.GSR = "ENABLED";
    FD1S3DX a_i3 (.D(a_31__N_2861[3]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i3.GSR = "ENABLED";
    FD1S3DX a_i4 (.D(a_31__N_2861[4]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i4.GSR = "ENABLED";
    FD1S3DX a_i5 (.D(a_31__N_2861[5]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i5.GSR = "ENABLED";
    FD1S3DX a_i6 (.D(a_31__N_2861[6]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i6.GSR = "ENABLED";
    FD1S3DX a_i7 (.D(a_31__N_2861[7]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i7.GSR = "ENABLED";
    FD1S3DX a_i8 (.D(a_31__N_2861[8]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i8.GSR = "ENABLED";
    FD1S3DX a_i9 (.D(a_31__N_2861[9]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i9.GSR = "ENABLED";
    FD1S3DX a_i10 (.D(a_31__N_2861[10]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i10.GSR = "ENABLED";
    FD1S3DX a_i11 (.D(a_31__N_2861[11]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i11.GSR = "ENABLED";
    FD1S3DX a_i12 (.D(a_31__N_2861[12]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i12.GSR = "ENABLED";
    FD1S3DX a_i13 (.D(a_31__N_2861[13]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i13.GSR = "ENABLED";
    FD1S3DX a_i14 (.D(a_31__N_2861[14]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i14.GSR = "ENABLED";
    FD1S3DX a_i15 (.D(a_31__N_2861[15]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i15.GSR = "ENABLED";
    FD1S3DX a_i16 (.D(a_31__N_2861[16]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i16.GSR = "ENABLED";
    FD1S3DX a_i17 (.D(a_31__N_2861[17]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i17.GSR = "ENABLED";
    FD1S3DX a_i18 (.D(a_31__N_2861[18]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i18.GSR = "ENABLED";
    FD1S3DX a_i19 (.D(a_31__N_2861[19]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i19.GSR = "ENABLED";
    FD1S3DX a_i20 (.D(a_31__N_2861[20]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i20.GSR = "ENABLED";
    FD1S3DX a_i21 (.D(a_31__N_2861[21]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i21.GSR = "ENABLED";
    FD1S3DX a_i22 (.D(a_31__N_2861[22]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i22.GSR = "ENABLED";
    FD1S3DX a_i23 (.D(a_31__N_2861[23]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i23.GSR = "ENABLED";
    FD1S3DX a_i24 (.D(a_31__N_2861[24]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i24.GSR = "ENABLED";
    FD1S3DX a_i25 (.D(a_31__N_2861[25]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i25.GSR = "ENABLED";
    FD1S3DX a_i26 (.D(a_31__N_2861[26]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i26.GSR = "ENABLED";
    FD1S3DX a_i27 (.D(a_31__N_2861[27]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i27.GSR = "ENABLED";
    FD1S3DX a_i28 (.D(a_31__N_2861[28]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i28.GSR = "ENABLED";
    FD1S3DX a_i29 (.D(a_31__N_2861[29]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i29.GSR = "ENABLED";
    FD1S3DX a_i30 (.D(a_31__N_2861[30]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(a[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i30.GSR = "ENABLED";
    FD1S3DX a_i31 (.D(a_31__N_2861[31]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\a[31] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i31.GSR = "ENABLED";
    FD1S3DX result_x_i1 (.D(result_x_31__N_2797[1]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i1.GSR = "ENABLED";
    FD1S3DX result_x_i2 (.D(result_x_31__N_2797[2]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i2.GSR = "ENABLED";
    FD1S3DX result_x_i3 (.D(result_x_31__N_2797[3]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i3.GSR = "ENABLED";
    FD1S3DX result_x_i4 (.D(result_x_31__N_2797[4]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i4.GSR = "ENABLED";
    FD1S3DX result_x_i5 (.D(result_x_31__N_2797[5]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i5.GSR = "ENABLED";
    FD1S3DX result_x_i6 (.D(result_x_31__N_2797[6]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i6.GSR = "ENABLED";
    FD1S3DX result_x_i7 (.D(result_x_31__N_2797[7]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i7.GSR = "ENABLED";
    FD1S3DX result_x_i8 (.D(result_x_31__N_2797[8]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i8.GSR = "ENABLED";
    FD1S3DX result_x_i9 (.D(result_x_31__N_2797[9]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i9.GSR = "ENABLED";
    FD1S3DX result_x_i10 (.D(result_x_31__N_2797[10]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i10.GSR = "ENABLED";
    FD1S3DX result_x_i11 (.D(result_x_31__N_2797[11]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i11.GSR = "ENABLED";
    FD1S3DX result_x_i12 (.D(result_x_31__N_2797[12]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i12.GSR = "ENABLED";
    FD1S3DX result_x_i13 (.D(result_x_31__N_2797[13]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i13.GSR = "ENABLED";
    FD1S3DX result_x_i14 (.D(result_x_31__N_2797[14]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i14.GSR = "ENABLED";
    FD1S3DX result_x_i15 (.D(result_x_31__N_2797[15]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i15.GSR = "ENABLED";
    FD1S3DX result_x_i16 (.D(result_x_31__N_2797[16]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i16.GSR = "ENABLED";
    FD1S3DX result_x_i17 (.D(result_x_31__N_2797[17]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i17.GSR = "ENABLED";
    FD1S3DX result_x_i18 (.D(result_x_31__N_2797[18]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i18.GSR = "ENABLED";
    FD1S3DX result_x_i19 (.D(result_x_31__N_2797[19]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i19.GSR = "ENABLED";
    FD1S3DX result_x_i20 (.D(result_x_31__N_2797[20]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i20.GSR = "ENABLED";
    FD1S3DX result_x_i21 (.D(result_x_31__N_2797[21]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i21.GSR = "ENABLED";
    FD1S3DX result_x_i22 (.D(result_x_31__N_2797[22]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i22.GSR = "ENABLED";
    FD1S3DX result_x_i23 (.D(result_x_31__N_2797[23]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i23.GSR = "ENABLED";
    FD1S3DX result_x_i24 (.D(result_x_31__N_2797[24]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i24.GSR = "ENABLED";
    FD1S3DX result_x_i25 (.D(result_x_31__N_2797[25]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i25.GSR = "ENABLED";
    FD1S3DX result_x_i26 (.D(result_x_31__N_2797[26]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i26.GSR = "ENABLED";
    FD1S3DX result_x_i27 (.D(result_x_31__N_2797[27]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i27.GSR = "ENABLED";
    FD1S3DX result_x_i28 (.D(result_x_31__N_2797[28]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i28.GSR = "ENABLED";
    FD1S3DX result_x_i29 (.D(result_x_31__N_2797[29]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i29.GSR = "ENABLED";
    FD1S3DX result_x_i30 (.D(result_x_31__N_2797[30]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i30.GSR = "ENABLED";
    FD1S3DX result_x_i31 (.D(result_x_31__N_2797[31]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(mc_result_x[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i31.GSR = "ENABLED";
    FD1S3DX cycles_i1 (.D(cycles_5__N_2928[1]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(cycles[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam cycles_i1.GSR = "ENABLED";
    FD1S3DX cycles_i2 (.D(cycles_5__N_2928[2]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(cycles[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam cycles_i2.GSR = "ENABLED";
    FD1S3DX cycles_i3 (.D(cycles_5__N_2928[3]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(cycles[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam cycles_i3.GSR = "ENABLED";
    FD1S3DX cycles_i4 (.D(cycles_5__N_2928[4]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(cycles[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam cycles_i4.GSR = "ENABLED";
    FD1S3DX cycles_i5 (.D(cycles_5__N_2928[5]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(cycles[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam cycles_i5.GSR = "ENABLED";
    CCU2C equal_30408_34 (.A0(n31889), .B0(n31888), .C0(n31887), .D0(n31886), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n35552), 
          .S1(divide_by_zero_x_N_3086));
    defparam equal_30408_34.INIT0 = 16'h8000;
    defparam equal_30408_34.INIT1 = 16'h0000;
    defparam equal_30408_34.INJECT1_0 = "YES";
    defparam equal_30408_34.INJECT1_1 = "NO";
    CCU2C equal_30408_33 (.A0(n31881), .B0(n31880), .C0(n31879), .D0(n31878), 
          .A1(n31885), .B1(n31884), .C1(n31883), .D1(n31882), .CIN(n35551), 
          .COUT(n35552));
    defparam equal_30408_33.INIT0 = 16'h8000;
    defparam equal_30408_33.INIT1 = 16'h8000;
    defparam equal_30408_33.INJECT1_0 = "YES";
    defparam equal_30408_33.INJECT1_1 = "YES";
    CCU2C equal_30408_31 (.A0(n31873), .B0(n31872), .C0(n31871), .D0(n31870), 
          .A1(n31877), .B1(n31876), .C1(n31875), .D1(n31874), .CIN(n35550), 
          .COUT(n35551));
    defparam equal_30408_31.INIT0 = 16'h8000;
    defparam equal_30408_31.INIT1 = 16'h8000;
    defparam equal_30408_31.INJECT1_0 = "YES";
    defparam equal_30408_31.INJECT1_1 = "YES";
    CCU2C equal_30408_29 (.A0(n31865), .B0(n31864), .C0(n31863), .D0(n31862), 
          .A1(n31869), .B1(n31868), .C1(n31867), .D1(n31866), .CIN(n35549), 
          .COUT(n35550));
    defparam equal_30408_29.INIT0 = 16'h8000;
    defparam equal_30408_29.INIT1 = 16'h8000;
    defparam equal_30408_29.INJECT1_0 = "YES";
    defparam equal_30408_29.INJECT1_1 = "YES";
    CCU2C equal_30408_0 (.A0(n31858), .B0(n41396), .C0(GND_net), .D0(VCC_net), 
          .A1(n31861), .B1(n31860), .C1(n31859), .D1(divide_by_zero_x_N_3090), 
          .COUT(n35549));
    defparam equal_30408_0.INIT0 = 16'h0008;
    defparam equal_30408_0.INIT1 = 16'h8000;
    defparam equal_30408_0.INJECT1_0 = "NO";
    defparam equal_30408_0.INJECT1_1 = "YES";
    LUT4 i4059_4_lut (.A(cycles_5__N_2936), .B(n32636), .C(divide_by_zero_x_N_3090), 
         .D(n15), .Z(n9349)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A ((D)+!B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i4059_4_lut.init = 16'h0ace;
    LUT4 divide_by_zero_x_I_126_4_lut (.A(n35380), .B(n41231), .C(cycles[0]), 
         .D(cycles[5]), .Z(divide_by_zero_x_N_3090)) /* synthesis lut_function=(A (B)+!A (B+!(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(244[17:69])
    defparam divide_by_zero_x_I_126_4_lut.init = 16'hcccd;
    LUT4 i1_4_lut (.A(cycles[3]), .B(cycles[2]), .C(cycles[4]), .D(cycles[1]), 
         .Z(n35380)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(244[17:48])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_991 (.A(state[0]), .B(cycles_5__N_2936), .Z(n41396)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_2_lut_rep_991.init = 16'heeee;
    LUT4 i4031_2_lut_3_lut (.A(state[0]), .B(cycles_5__N_2936), .C(divide_by_zero_x_N_3090), 
         .Z(n9312)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i4031_2_lut_3_lut.init = 16'he0e0;
    LUT4 select_1205_Select_1_i1_3_lut_4_lut (.A(state[0]), .B(cycles_5__N_2936), 
         .C(cycles[0]), .D(cycles[1]), .Z(n1_adj_6104)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1205_Select_1_i1_3_lut_4_lut.init = 16'he00e;
    LUT4 select_1205_Select_2_i1_3_lut_4_lut (.A(state[0]), .B(cycles_5__N_2936), 
         .C(n41445), .D(cycles[2]), .Z(n1_adj_6105)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1205_Select_2_i1_3_lut_4_lut.init = 16'he00e;
    LUT4 select_1202_Select_1_i3_4_lut (.A(n1_adj_6106), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[1]), .Z(p_31__N_2829[1])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_1_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_1_i1_4_lut (.A(t[1]), .B(n41396), .C(p[0]), 
         .D(t[32]), .Z(n1_adj_6106)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_1_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_2_i3_4_lut (.A(n1_adj_6107), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[2]), .Z(p_31__N_2829[2])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_2_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_2_i1_4_lut (.A(t[2]), .B(n41396), .C(p[1]), 
         .D(t[32]), .Z(n1_adj_6107)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_2_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_3_i3_4_lut (.A(n1_adj_6108), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[3]), .Z(p_31__N_2829[3])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_3_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_3_i1_4_lut (.A(t[3]), .B(n41396), .C(p[2]), 
         .D(t[32]), .Z(n1_adj_6108)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_3_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_4_i3_4_lut (.A(n1_adj_6109), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[4]), .Z(p_31__N_2829[4])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_4_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_4_i1_4_lut (.A(t[4]), .B(n41396), .C(p[3]), 
         .D(t[32]), .Z(n1_adj_6109)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_4_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_5_i3_4_lut (.A(n1_adj_6110), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[5]), .Z(p_31__N_2829[5])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_5_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_5_i1_4_lut (.A(t[5]), .B(n41396), .C(p[4]), 
         .D(t[32]), .Z(n1_adj_6110)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_5_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_6_i3_4_lut (.A(n1_adj_6111), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[6]), .Z(p_31__N_2829[6])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_6_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_6_i1_4_lut (.A(t[6]), .B(n41396), .C(p[5]), 
         .D(t[32]), .Z(n1_adj_6111)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_6_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_7_i3_4_lut (.A(n1_adj_6112), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[7]), .Z(p_31__N_2829[7])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_7_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_7_i1_4_lut (.A(t[7]), .B(n41396), .C(p[6]), 
         .D(t[32]), .Z(n1_adj_6112)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_7_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_8_i3_4_lut (.A(n1_adj_6113), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[8]), .Z(p_31__N_2829[8])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_8_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_8_i1_4_lut (.A(t[8]), .B(n41396), .C(p[7]), 
         .D(t[32]), .Z(n1_adj_6113)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_8_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_9_i3_4_lut (.A(n1_adj_6114), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[9]), .Z(p_31__N_2829[9])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_9_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_9_i1_4_lut (.A(t[9]), .B(n41396), .C(p[8]), 
         .D(t[32]), .Z(n1_adj_6114)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_9_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_10_i3_4_lut (.A(n1_adj_6115), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[10]), .Z(p_31__N_2829[10])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_10_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_10_i1_4_lut (.A(t[10]), .B(n41396), .C(p[9]), 
         .D(t[32]), .Z(n1_adj_6115)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_10_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_11_i3_4_lut (.A(n1_adj_6116), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[11]), .Z(p_31__N_2829[11])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_11_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_11_i1_4_lut (.A(t[11]), .B(n41396), .C(p[10]), 
         .D(t[32]), .Z(n1_adj_6116)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_11_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_12_i3_4_lut (.A(n1_adj_6117), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[12]), .Z(p_31__N_2829[12])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_12_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_12_i1_4_lut (.A(t[12]), .B(n41396), .C(p[11]), 
         .D(t[32]), .Z(n1_adj_6117)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_12_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_13_i3_4_lut (.A(n1_adj_6118), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[13]), .Z(p_31__N_2829[13])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_13_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_13_i1_4_lut (.A(t[13]), .B(n41396), .C(p[12]), 
         .D(t[32]), .Z(n1_adj_6118)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_13_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_14_i3_4_lut (.A(n1_adj_6119), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[14]), .Z(p_31__N_2829[14])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_14_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_14_i1_4_lut (.A(t[14]), .B(n41396), .C(p[13]), 
         .D(t[32]), .Z(n1_adj_6119)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_14_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_15_i3_4_lut (.A(n1_adj_6120), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[15]), .Z(p_31__N_2829[15])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_15_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_15_i1_4_lut (.A(t[15]), .B(n41396), .C(p[14]), 
         .D(t[32]), .Z(n1_adj_6120)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_15_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_16_i3_4_lut (.A(n1_adj_6121), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[16]), .Z(p_31__N_2829[16])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_16_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_16_i1_4_lut (.A(t[16]), .B(n41396), .C(p[15]), 
         .D(t[32]), .Z(n1_adj_6121)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_16_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_17_i3_4_lut (.A(n1_adj_6122), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[17]), .Z(p_31__N_2829[17])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_17_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_17_i1_4_lut (.A(t[17]), .B(n41396), .C(p[16]), 
         .D(t[32]), .Z(n1_adj_6122)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_17_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_18_i3_4_lut (.A(n1_adj_6123), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[18]), .Z(p_31__N_2829[18])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_18_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_18_i1_4_lut (.A(t[18]), .B(n41396), .C(p[17]), 
         .D(t[32]), .Z(n1_adj_6123)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_18_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_19_i3_4_lut (.A(n1_adj_6124), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[19]), .Z(p_31__N_2829[19])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_19_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_19_i1_4_lut (.A(t[19]), .B(n41396), .C(p[18]), 
         .D(t[32]), .Z(n1_adj_6124)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_19_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_20_i3_4_lut (.A(n1_adj_6125), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[20]), .Z(p_31__N_2829[20])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_20_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_20_i1_4_lut (.A(t[20]), .B(n41396), .C(p[19]), 
         .D(t[32]), .Z(n1_adj_6125)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_20_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_21_i3_4_lut (.A(n1_adj_6126), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[21]), .Z(p_31__N_2829[21])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_21_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_21_i1_4_lut (.A(t[21]), .B(n41396), .C(p[20]), 
         .D(t[32]), .Z(n1_adj_6126)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_21_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_22_i3_4_lut (.A(n1_adj_6127), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[22]), .Z(p_31__N_2829[22])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_22_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_22_i1_4_lut (.A(t[22]), .B(n41396), .C(p[21]), 
         .D(t[32]), .Z(n1_adj_6127)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_22_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_23_i3_4_lut (.A(n1_adj_6128), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[23]), .Z(p_31__N_2829[23])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_23_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_23_i1_4_lut (.A(t[23]), .B(n41396), .C(p[22]), 
         .D(t[32]), .Z(n1_adj_6128)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_23_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_24_i3_4_lut (.A(n1_adj_6129), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[24]), .Z(p_31__N_2829[24])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_24_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_24_i1_4_lut (.A(t[24]), .B(n41396), .C(p[23]), 
         .D(t[32]), .Z(n1_adj_6129)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_24_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_25_i3_4_lut (.A(n1_adj_6130), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[25]), .Z(p_31__N_2829[25])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_25_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_25_i1_4_lut (.A(t[25]), .B(n41396), .C(p[24]), 
         .D(t[32]), .Z(n1_adj_6130)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_25_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_26_i3_4_lut (.A(n1_adj_6131), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[26]), .Z(p_31__N_2829[26])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_26_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_26_i1_4_lut (.A(t[26]), .B(n41396), .C(p[25]), 
         .D(t[32]), .Z(n1_adj_6131)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_26_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_27_i3_4_lut (.A(n1_adj_6132), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[27]), .Z(p_31__N_2829[27])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_27_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_27_i1_4_lut (.A(t[27]), .B(n41396), .C(p[26]), 
         .D(t[32]), .Z(n1_adj_6132)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_27_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_28_i3_4_lut (.A(n1_adj_6133), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[28]), .Z(p_31__N_2829[28])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_28_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_28_i1_4_lut (.A(t[28]), .B(n41396), .C(p[27]), 
         .D(t[32]), .Z(n1_adj_6133)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_28_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_29_i3_4_lut (.A(n1_adj_6134), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[29]), .Z(p_31__N_2829[29])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_29_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_29_i1_4_lut (.A(t[29]), .B(n41396), .C(p[28]), 
         .D(t[32]), .Z(n1_adj_6134)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_29_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_30_i3_4_lut (.A(n1_adj_6135), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[30]), .Z(p_31__N_2829[30])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_30_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_30_i1_4_lut (.A(t[30]), .B(n41396), .C(p[29]), 
         .D(t[32]), .Z(n1_adj_6135)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_30_i1_4_lut.init = 16'hc088;
    LUT4 select_1202_Select_31_i3_4_lut (.A(n1_adj_6136), .B(cycles_5__N_2934), 
         .C(n45183), .D(p_c[31]), .Z(p_31__N_2829[31])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_31_i3_4_lut.init = 16'heaaa;
    LUT4 select_1202_Select_31_i1_4_lut (.A(t[31]), .B(n41396), .C(p[30]), 
         .D(t[32]), .Z(n1_adj_6136)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_31_i1_4_lut.init = 16'hc088;
    LUT4 i2_4_lut (.A(a_31__N_3014[1]), .B(a[0]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[1])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut.init = 16'heca0;
    LUT4 mux_13_i2_3_lut (.A(d_result_0[1]), .B(a[1]), .C(n45183), .Z(a_31__N_3014[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_511 (.A(a[1]), .B(a_31__N_3014[2]), .C(n41396), 
         .D(cycles_5__N_2934), .Z(a_31__N_2861[2])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_511.init = 16'heca0;
    LUT4 mux_13_i3_3_lut (.A(d_result_0[2]), .B(a[2]), .C(n45183), .Z(a_31__N_3014[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i3_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_512 (.A(a_31__N_3014[3]), .B(a[2]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[3])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_512.init = 16'heca0;
    LUT4 mux_13_i4_3_lut (.A(d_result_0[3]), .B(a[3]), .C(n45183), .Z(a_31__N_3014[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i4_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_513 (.A(a_31__N_3014[4]), .B(a[3]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[4])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_513.init = 16'heca0;
    LUT4 mux_13_i5_3_lut (.A(d_result_0[4]), .B(a[4]), .C(n45183), .Z(a_31__N_3014[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i5_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_514 (.A(a_31__N_3014[5]), .B(a[4]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[5])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_514.init = 16'heca0;
    LUT4 mux_13_i6_3_lut (.A(d_result_0[5]), .B(a[5]), .C(n45183), .Z(a_31__N_3014[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i6_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_515 (.A(a[5]), .B(a_31__N_3014[6]), .C(n41396), 
         .D(cycles_5__N_2934), .Z(a_31__N_2861[6])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_515.init = 16'heca0;
    LUT4 mux_13_i7_3_lut (.A(d_result_0[6]), .B(a[6]), .C(n45183), .Z(a_31__N_3014[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i7_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_516 (.A(a_31__N_3014[7]), .B(a[6]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[7])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_516.init = 16'heca0;
    LUT4 mux_13_i8_3_lut (.A(d_result_0[7]), .B(a[7]), .C(n45183), .Z(a_31__N_3014[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i8_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_517 (.A(a_31__N_3014[8]), .B(a[7]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[8])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_517.init = 16'heca0;
    LUT4 mux_13_i9_3_lut (.A(d_result_0[8]), .B(a[8]), .C(n45183), .Z(a_31__N_3014[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i9_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_518 (.A(a[8]), .B(a_31__N_3014[9]), .C(n41396), 
         .D(cycles_5__N_2934), .Z(a_31__N_2861[9])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_518.init = 16'heca0;
    LUT4 mux_13_i10_3_lut (.A(d_result_0[9]), .B(a[9]), .C(n45183), .Z(a_31__N_3014[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i10_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_519 (.A(a_31__N_3014[10]), .B(a[9]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[10])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_519.init = 16'heca0;
    LUT4 mux_13_i11_3_lut (.A(d_result_0[10]), .B(a[10]), .C(n45183), 
         .Z(a_31__N_3014[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i11_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_520 (.A(a_31__N_3014[11]), .B(a[10]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[11])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_520.init = 16'heca0;
    LUT4 mux_13_i12_3_lut (.A(d_result_0[11]), .B(a[11]), .C(n45183), 
         .Z(a_31__N_3014[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i12_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_521 (.A(a[11]), .B(a_31__N_3014[12]), .C(n41396), 
         .D(cycles_5__N_2934), .Z(a_31__N_2861[12])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_521.init = 16'heca0;
    LUT4 mux_13_i13_3_lut (.A(d_result_0[12]), .B(a[12]), .C(n45183), 
         .Z(a_31__N_3014[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i13_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_522 (.A(a_31__N_3014[13]), .B(a[12]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[13])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_522.init = 16'heca0;
    LUT4 mux_13_i14_3_lut (.A(d_result_0[13]), .B(a[13]), .C(n45183), 
         .Z(a_31__N_3014[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i14_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_523 (.A(a[13]), .B(a_31__N_3014[14]), .C(n41396), 
         .D(cycles_5__N_2934), .Z(a_31__N_2861[14])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_523.init = 16'heca0;
    LUT4 mux_13_i15_3_lut (.A(d_result_0[14]), .B(a[14]), .C(n45183), 
         .Z(a_31__N_3014[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i15_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_524 (.A(a[14]), .B(a_31__N_3014[15]), .C(n41396), 
         .D(cycles_5__N_2934), .Z(a_31__N_2861[15])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_524.init = 16'heca0;
    LUT4 mux_13_i16_3_lut (.A(d_result_0[15]), .B(a[15]), .C(n45183), 
         .Z(a_31__N_3014[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i16_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_525 (.A(a_31__N_3014[16]), .B(a[15]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[16])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_525.init = 16'heca0;
    LUT4 mux_13_i17_3_lut (.A(d_result_0[16]), .B(a[16]), .C(n45183), 
         .Z(a_31__N_3014[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i17_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_526 (.A(a[16]), .B(a_31__N_3014[17]), .C(n41396), 
         .D(cycles_5__N_2934), .Z(a_31__N_2861[17])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_526.init = 16'heca0;
    LUT4 mux_13_i18_3_lut (.A(d_result_0[17]), .B(a[17]), .C(n45183), 
         .Z(a_31__N_3014[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i18_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_527 (.A(a_31__N_3014[18]), .B(a[17]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[18])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_527.init = 16'heca0;
    LUT4 mux_13_i19_3_lut (.A(d_result_0[18]), .B(a[18]), .C(n45183), 
         .Z(a_31__N_3014[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i19_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_528 (.A(a_31__N_3014[19]), .B(a[18]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[19])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_528.init = 16'heca0;
    LUT4 mux_13_i20_3_lut (.A(d_result_0[19]), .B(a[19]), .C(n45183), 
         .Z(a_31__N_3014[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i20_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_529 (.A(a[19]), .B(a_31__N_3014[20]), .C(n41396), 
         .D(cycles_5__N_2934), .Z(a_31__N_2861[20])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_529.init = 16'heca0;
    LUT4 select_1202_Select_0_i3_4_lut (.A(n1_adj_6137), .B(cycles_5__N_2934), 
         .C(n45183), .D(p[0]), .Z(p_31__N_2829[0])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_0_i3_4_lut.init = 16'heaaa;
    LUT4 mux_13_i21_3_lut (.A(d_result_0[20]), .B(a[20]), .C(n45183), 
         .Z(a_31__N_3014[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i21_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_530 (.A(a_31__N_3014[21]), .B(a[20]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[21])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_530.init = 16'heca0;
    LUT4 mux_13_i22_3_lut (.A(d_result_0[21]), .B(a[21]), .C(n45183), 
         .Z(a_31__N_3014[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i22_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_531 (.A(a_31__N_3014[22]), .B(a[21]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[22])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_531.init = 16'heca0;
    LUT4 select_1202_Select_0_i1_4_lut (.A(t[0]), .B(n41396), .C(\a[31] ), 
         .D(t[32]), .Z(n1_adj_6137)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1202_Select_0_i1_4_lut.init = 16'hc088;
    LUT4 mux_13_i23_3_lut (.A(d_result_0[22]), .B(a[22]), .C(n45183), 
         .Z(a_31__N_3014[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i23_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_532 (.A(a_31__N_3014[23]), .B(a[22]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[23])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_532.init = 16'heca0;
    LUT4 i1_4_lut_adj_533 (.A(a_31__N_3014[0]), .B(t[32]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[0])) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A !(B+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_533.init = 16'hb3a0;
    LUT4 mux_13_i24_3_lut (.A(d_result_0[23]), .B(a[23]), .C(n45183), 
         .Z(a_31__N_3014[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i24_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_534 (.A(a_31__N_3014[24]), .B(a[23]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[24])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_534.init = 16'heca0;
    LUT4 mux_13_i25_3_lut (.A(d_result_0[24]), .B(a[24]), .C(n45183), 
         .Z(a_31__N_3014[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i25_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_535 (.A(a_31__N_3014[25]), .B(a[24]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[25])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_535.init = 16'heca0;
    LUT4 mux_13_i26_3_lut (.A(d_result_0[25]), .B(a[25]), .C(n45183), 
         .Z(a_31__N_3014[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i26_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_536 (.A(a[25]), .B(a_31__N_3014[26]), .C(n41396), 
         .D(cycles_5__N_2934), .Z(a_31__N_2861[26])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_536.init = 16'heca0;
    LUT4 mux_13_i27_3_lut (.A(d_result_0[26]), .B(a[26]), .C(n45183), 
         .Z(a_31__N_3014[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i27_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_537 (.A(a[26]), .B(a_31__N_3014[27]), .C(n41396), 
         .D(cycles_5__N_2934), .Z(a_31__N_2861[27])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_537.init = 16'heca0;
    LUT4 mux_13_i1_3_lut (.A(d_result_0[0]), .B(a[0]), .C(n45183), .Z(a_31__N_3014[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i1_3_lut.init = 16'hcaca;
    LUT4 mux_13_i28_3_lut (.A(d_result_0[27]), .B(a[27]), .C(n45183), 
         .Z(a_31__N_3014[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i28_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_538 (.A(a_31__N_3014[28]), .B(a[27]), .C(cycles_5__N_2934), 
         .D(n41396), .Z(a_31__N_2861[28])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_538.init = 16'heca0;
    LUT4 i2_4_lut_adj_539 (.A(n1_adj_6138), .B(mc_result_x[0]), .C(n2), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[0])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_539.init = 16'hfefa;
    LUT4 mux_13_i29_3_lut (.A(d_result_0[28]), .B(a[28]), .C(n45183), 
         .Z(a_31__N_3014[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i29_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_540 (.A(a[28]), .B(a_31__N_3014[29]), .C(n41396), 
         .D(cycles_5__N_2934), .Z(a_31__N_2861[29])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_540.init = 16'heca0;
    LUT4 mux_13_i30_3_lut (.A(d_result_0[29]), .B(a[29]), .C(n45183), 
         .Z(a_31__N_3014[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i30_3_lut.init = 16'hcaca;
    LUT4 select_519_Select_0_i1_2_lut (.A(p[0]), .B(cycles_5__N_2936), .Z(n1_adj_6138)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_0_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_0_i2_2_lut (.A(a[0]), .B(state[0]), .Z(n2)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_0_i2_2_lut.init = 16'h8888;
    LUT4 i11_4_lut (.A(n41396), .B(n45183), .C(cycles[0]), .D(cycles_5__N_2934), 
         .Z(cycles_5__N_2928[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i11_4_lut.init = 16'hca0a;
    LUT4 i1_4_lut_adj_541 (.A(a[29]), .B(a_31__N_3014[30]), .C(n41396), 
         .D(cycles_5__N_2934), .Z(a_31__N_2861[30])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_541.init = 16'heca0;
    LUT4 mux_13_i31_3_lut (.A(d_result_0[30]), .B(a[30]), .C(n45183), 
         .Z(a_31__N_3014[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i31_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_542 (.A(a[30]), .B(a_31__N_3014[31]), .C(n41396), 
         .D(cycles_5__N_2934), .Z(a_31__N_2861[31])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_542.init = 16'heca0;
    LUT4 mux_13_i32_3_lut (.A(d_result_0[31]), .B(\a[31] ), .C(n45183), 
         .Z(a_31__N_3014[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(194[13] 228[16])
    defparam mux_13_i32_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut (.A(mc_result_x[1]), .B(n4), .C(cycles_5__N_2934), .Z(result_x_31__N_2797[1])) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_543 (.A(a[1]), .B(p[1]), .C(state[0]), .D(cycles_5__N_2936), 
         .Z(n4)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_543.init = 16'heca0;
    LUT4 i2_4_lut_adj_544 (.A(n1_adj_6139), .B(mc_result_x[2]), .C(n2_adj_6140), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[2])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_544.init = 16'hfefa;
    LUT4 select_519_Select_2_i1_2_lut (.A(p[2]), .B(cycles_5__N_2936), .Z(n1_adj_6139)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_2_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_2_i2_2_lut (.A(a[2]), .B(state[0]), .Z(n2_adj_6140)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_2_i2_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_545 (.A(n1_adj_6141), .B(n2_adj_6142), .C(mc_result_x[3]), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[3])) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_545.init = 16'hfeee;
    LUT4 select_519_Select_3_i1_2_lut (.A(p[3]), .B(cycles_5__N_2936), .Z(n1_adj_6141)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_3_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_3_i2_2_lut (.A(a[3]), .B(state[0]), .Z(n2_adj_6142)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_3_i2_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_546 (.A(n1_adj_6143), .B(mc_result_x[4]), .C(n2_adj_6144), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[4])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_546.init = 16'hfefa;
    LUT4 select_519_Select_4_i1_2_lut (.A(p[4]), .B(cycles_5__N_2936), .Z(n1_adj_6143)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_4_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_4_i2_2_lut (.A(a[4]), .B(state[0]), .Z(n2_adj_6144)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_4_i2_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_547 (.A(n1_adj_6145), .B(n2_adj_6146), .C(mc_result_x[5]), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[5])) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_547.init = 16'hfeee;
    LUT4 select_519_Select_5_i1_2_lut (.A(p[5]), .B(cycles_5__N_2936), .Z(n1_adj_6145)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_5_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_5_i2_2_lut (.A(a[5]), .B(state[0]), .Z(n2_adj_6146)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_5_i2_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_548 (.A(n1_adj_6147), .B(mc_result_x[6]), .C(n2_adj_6148), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[6])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_548.init = 16'hfefa;
    LUT4 select_519_Select_6_i1_2_lut (.A(p[6]), .B(cycles_5__N_2936), .Z(n1_adj_6147)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_6_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_6_i2_2_lut (.A(a[6]), .B(state[0]), .Z(n2_adj_6148)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_6_i2_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_549 (.A(n1_adj_6149), .B(mc_result_x[7]), .C(n2_adj_6150), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[7])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_549.init = 16'hfefa;
    LUT4 select_519_Select_7_i1_2_lut (.A(p[7]), .B(cycles_5__N_2936), .Z(n1_adj_6149)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_7_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_7_i2_2_lut (.A(a[7]), .B(state[0]), .Z(n2_adj_6150)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_7_i2_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_550 (.A(n1_adj_6151), .B(mc_result_x[8]), .C(n2_adj_6152), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[8])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_550.init = 16'hfefa;
    LUT4 select_519_Select_8_i1_2_lut (.A(p[8]), .B(cycles_5__N_2936), .Z(n1_adj_6151)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_8_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_8_i2_2_lut (.A(a[8]), .B(state[0]), .Z(n2_adj_6152)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_8_i2_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_551 (.A(n1_adj_6153), .B(n2_adj_6154), .C(mc_result_x[9]), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[9])) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_551.init = 16'hfeee;
    LUT4 select_519_Select_9_i1_2_lut (.A(p[9]), .B(cycles_5__N_2936), .Z(n1_adj_6153)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_9_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_9_i2_2_lut (.A(a[9]), .B(state[0]), .Z(n2_adj_6154)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_9_i2_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_552 (.A(n1_adj_6155), .B(mc_result_x[10]), .C(n2_adj_6156), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[10])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_552.init = 16'hfefa;
    LUT4 select_519_Select_10_i1_2_lut (.A(p[10]), .B(cycles_5__N_2936), 
         .Z(n1_adj_6155)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_10_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_10_i2_2_lut (.A(a[10]), .B(state[0]), .Z(n2_adj_6156)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_10_i2_2_lut.init = 16'h8888;
    LUT4 i2_3_lut_adj_553 (.A(mc_result_x[11]), .B(n4_adj_6157), .C(cycles_5__N_2934), 
         .Z(result_x_31__N_2797[11])) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_3_lut_adj_553.init = 16'hecec;
    LUT4 i1_4_lut_adj_554 (.A(a[11]), .B(p[11]), .C(state[0]), .D(cycles_5__N_2936), 
         .Z(n4_adj_6157)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_554.init = 16'heca0;
    LUT4 i2_4_lut_adj_555 (.A(n1_adj_6158), .B(n2_adj_6159), .C(mc_result_x[12]), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[12])) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_555.init = 16'hfeee;
    LUT4 select_519_Select_12_i1_2_lut (.A(p[12]), .B(cycles_5__N_2936), 
         .Z(n1_adj_6158)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_12_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_12_i2_2_lut (.A(a[12]), .B(state[0]), .Z(n2_adj_6159)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_12_i2_2_lut.init = 16'h8888;
    LUT4 i2_3_lut_adj_556 (.A(mc_result_x[13]), .B(n4_adj_6160), .C(cycles_5__N_2934), 
         .Z(result_x_31__N_2797[13])) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_3_lut_adj_556.init = 16'hecec;
    LUT4 i1_4_lut_adj_557 (.A(a[13]), .B(p[13]), .C(state[0]), .D(cycles_5__N_2936), 
         .Z(n4_adj_6160)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_557.init = 16'heca0;
    LUT4 i2_4_lut_adj_558 (.A(n1_adj_6161), .B(n2_adj_6162), .C(mc_result_x[14]), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[14])) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_558.init = 16'hfeee;
    LUT4 select_519_Select_14_i1_2_lut (.A(p[14]), .B(cycles_5__N_2936), 
         .Z(n1_adj_6161)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_14_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_14_i2_2_lut (.A(a[14]), .B(state[0]), .Z(n2_adj_6162)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_14_i2_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_559 (.A(n1_adj_6163), .B(mc_result_x[15]), .C(n2_adj_6164), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[15])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_559.init = 16'hfefa;
    LUT4 select_519_Select_15_i1_2_lut (.A(p[15]), .B(cycles_5__N_2936), 
         .Z(n1_adj_6163)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_15_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_15_i2_2_lut (.A(a[15]), .B(state[0]), .Z(n2_adj_6164)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_15_i2_2_lut.init = 16'h8888;
    LUT4 i2_3_lut_adj_560 (.A(mc_result_x[16]), .B(n4_adj_6165), .C(cycles_5__N_2934), 
         .Z(result_x_31__N_2797[16])) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_3_lut_adj_560.init = 16'hecec;
    LUT4 i1_4_lut_adj_561 (.A(a[16]), .B(p[16]), .C(state[0]), .D(cycles_5__N_2936), 
         .Z(n4_adj_6165)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_561.init = 16'heca0;
    LUT4 i2_4_lut_adj_562 (.A(n1_adj_6166), .B(mc_result_x[17]), .C(n2_adj_6167), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[17])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_562.init = 16'hfefa;
    LUT4 select_519_Select_17_i1_2_lut (.A(p[17]), .B(cycles_5__N_2936), 
         .Z(n1_adj_6166)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_17_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_17_i2_2_lut (.A(a[17]), .B(state[0]), .Z(n2_adj_6167)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_17_i2_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_563 (.A(n1_adj_6168), .B(mc_result_x[18]), .C(n2_adj_6169), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[18])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_563.init = 16'hfefa;
    LUT4 select_519_Select_18_i1_2_lut (.A(p[18]), .B(cycles_5__N_2936), 
         .Z(n1_adj_6168)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_18_i1_2_lut.init = 16'h8888;
    LUT4 select_518_Select_19_i2_2_lut (.A(a[18]), .B(state[0]), .Z(n2_adj_6169)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_518_Select_19_i2_2_lut.init = 16'h8888;
    LUT4 i2_3_lut_adj_564 (.A(mc_result_x[19]), .B(n4_adj_6170), .C(cycles_5__N_2934), 
         .Z(result_x_31__N_2797[19])) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_3_lut_adj_564.init = 16'hecec;
    LUT4 i1_4_lut_adj_565 (.A(a[19]), .B(p[19]), .C(state[0]), .D(cycles_5__N_2936), 
         .Z(n4_adj_6170)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_565.init = 16'heca0;
    LUT4 i2_4_lut_adj_566 (.A(n1_adj_6171), .B(mc_result_x[20]), .C(n2_adj_6172), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[20])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_566.init = 16'hfefa;
    LUT4 select_519_Select_20_i1_2_lut (.A(p[20]), .B(cycles_5__N_2936), 
         .Z(n1_adj_6171)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_20_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_20_i2_2_lut (.A(a[20]), .B(state[0]), .Z(n2_adj_6172)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_20_i2_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_567 (.A(n1_adj_6173), .B(n2_adj_6174), .C(mc_result_x[21]), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[21])) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_567.init = 16'hfeee;
    LUT4 select_519_Select_21_i1_2_lut (.A(p[21]), .B(cycles_5__N_2936), 
         .Z(n1_adj_6173)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_21_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_21_i2_2_lut (.A(a[21]), .B(state[0]), .Z(n2_adj_6174)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_21_i2_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_568 (.A(n1_adj_6175), .B(mc_result_x[22]), .C(n2_adj_6176), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[22])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_568.init = 16'hfefa;
    LUT4 select_519_Select_22_i1_2_lut (.A(p[22]), .B(cycles_5__N_2936), 
         .Z(n1_adj_6175)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_22_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_22_i2_2_lut (.A(a[22]), .B(state[0]), .Z(n2_adj_6176)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_22_i2_2_lut.init = 16'h8888;
    LUT4 i2_3_lut_adj_569 (.A(mc_result_x[23]), .B(n4_adj_6177), .C(cycles_5__N_2934), 
         .Z(result_x_31__N_2797[23])) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_3_lut_adj_569.init = 16'hecec;
    LUT4 i1_4_lut_adj_570 (.A(a[23]), .B(p[23]), .C(state[0]), .D(cycles_5__N_2936), 
         .Z(n4_adj_6177)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_570.init = 16'heca0;
    LUT4 i2_4_lut_adj_571 (.A(n1_adj_6178), .B(n2_adj_6179), .C(mc_result_x[24]), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[24])) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_571.init = 16'hfeee;
    LUT4 select_519_Select_24_i1_2_lut (.A(p[24]), .B(cycles_5__N_2936), 
         .Z(n1_adj_6178)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_24_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_24_i2_2_lut (.A(a[24]), .B(state[0]), .Z(n2_adj_6179)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_24_i2_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_572 (.A(n1_adj_6180), .B(n2_adj_6181), .C(mc_result_x[25]), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[25])) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_572.init = 16'hfeee;
    LUT4 select_519_Select_25_i1_2_lut (.A(p[25]), .B(cycles_5__N_2936), 
         .Z(n1_adj_6180)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_25_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_25_i2_2_lut (.A(a[25]), .B(state[0]), .Z(n2_adj_6181)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_25_i2_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_573 (.A(n1_adj_6182), .B(n2_adj_6183), .C(mc_result_x[26]), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[26])) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_573.init = 16'hfeee;
    LUT4 select_519_Select_26_i1_2_lut (.A(p[26]), .B(cycles_5__N_2936), 
         .Z(n1_adj_6182)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_26_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_26_i2_2_lut (.A(a[26]), .B(state[0]), .Z(n2_adj_6183)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_26_i2_2_lut.init = 16'h8888;
    LUT4 i2_3_lut_adj_574 (.A(mc_result_x[27]), .B(n4_adj_6184), .C(cycles_5__N_2934), 
         .Z(result_x_31__N_2797[27])) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_3_lut_adj_574.init = 16'hecec;
    LUT4 i1_4_lut_adj_575 (.A(a[27]), .B(p[27]), .C(state[0]), .D(cycles_5__N_2936), 
         .Z(n4_adj_6184)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_575.init = 16'heca0;
    LUT4 i2_3_lut_adj_576 (.A(mc_result_x[28]), .B(n4_adj_6185), .C(cycles_5__N_2934), 
         .Z(result_x_31__N_2797[28])) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_3_lut_adj_576.init = 16'hecec;
    LUT4 i1_4_lut_adj_577 (.A(a[28]), .B(p[28]), .C(state[0]), .D(cycles_5__N_2936), 
         .Z(n4_adj_6185)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_577.init = 16'heca0;
    LUT4 i2_3_lut_adj_578 (.A(mc_result_x[29]), .B(n4_adj_6186), .C(cycles_5__N_2934), 
         .Z(result_x_31__N_2797[29])) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_3_lut_adj_578.init = 16'hecec;
    LUT4 i1_4_lut_adj_579 (.A(a[29]), .B(p[29]), .C(state[0]), .D(cycles_5__N_2936), 
         .Z(n4_adj_6186)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i1_4_lut_adj_579.init = 16'heca0;
    LUT4 i2_4_lut_adj_580 (.A(n1_adj_6187), .B(mc_result_x[30]), .C(n2_adj_6188), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[30])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_580.init = 16'hfefa;
    LUT4 select_519_Select_30_i1_2_lut (.A(p[30]), .B(cycles_5__N_2936), 
         .Z(n1_adj_6187)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_30_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_30_i2_2_lut (.A(a[30]), .B(state[0]), .Z(n2_adj_6188)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_30_i2_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_581 (.A(n1_adj_6189), .B(n2_adj_6190), .C(mc_result_x[31]), 
         .D(cycles_5__N_2934), .Z(result_x_31__N_2797[31])) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i2_4_lut_adj_581.init = 16'hfeee;
    LUT4 select_519_Select_31_i1_2_lut (.A(p_c[31]), .B(cycles_5__N_2936), 
         .Z(n1_adj_6189)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_31_i1_2_lut.init = 16'h8888;
    LUT4 select_519_Select_31_i2_2_lut (.A(\a[31] ), .B(state[0]), .Z(n2_adj_6190)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_519_Select_31_i2_2_lut.init = 16'h8888;
    LUT4 select_1205_Select_1_i3_4_lut (.A(n1_adj_6104), .B(cycles_5__N_2934), 
         .C(n45183), .D(cycles[1]), .Z(cycles_5__N_2928[1])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1205_Select_1_i3_4_lut.init = 16'heaaa;
    LUT4 select_1205_Select_2_i3_4_lut (.A(n1_adj_6105), .B(cycles_5__N_2934), 
         .C(n45183), .D(cycles[2]), .Z(cycles_5__N_2928[2])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1205_Select_2_i3_4_lut.init = 16'heaaa;
    LUT4 select_1205_Select_3_i3_4_lut (.A(n1), .B(cycles_5__N_2934), .C(n45183), 
         .D(cycles[3]), .Z(cycles_5__N_2928[3])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1205_Select_3_i3_4_lut.init = 16'heaaa;
    LUT4 select_1205_Select_4_i3_4_lut (.A(n1_adj_6191), .B(cycles_5__N_2934), 
         .C(n45183), .D(cycles[4]), .Z(cycles_5__N_2928[4])) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1205_Select_4_i3_4_lut.init = 16'heaaa;
    LUT4 select_1205_Select_5_i3_4_lut (.A(n1_adj_6192), .B(cycles[5]), 
         .C(cycles_5__N_2934), .D(n45181), .Z(cycles_5__N_2928[5])) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1205_Select_5_i3_4_lut.init = 16'hfaea;
    LUT4 select_1205_Select_5_i1_4_lut (.A(cycles[5]), .B(n41396), .C(cycles[4]), 
         .D(n41293), .Z(n1_adj_6192)) /* synthesis lut_function=(A (B (C+(D)))+!A !((C+(D))+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam select_1205_Select_5_i1_4_lut.init = 16'h8884;
    LUT4 i26750_1_lut (.A(b[28]), .Z(n31889)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26750_1_lut.init = 16'h5555;
    LUT4 i26749_1_lut (.A(b[31]), .Z(n31888)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26749_1_lut.init = 16'h5555;
    LUT4 i26748_1_lut (.A(b[13]), .Z(n31887)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26748_1_lut.init = 16'h5555;
    LUT4 i26747_1_lut (.A(b[23]), .Z(n31886)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26747_1_lut.init = 16'h5555;
    LUT4 i26742_1_lut (.A(b[14]), .Z(n31881)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26742_1_lut.init = 16'h5555;
    LUT4 i26741_1_lut (.A(b[30]), .Z(n31880)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26741_1_lut.init = 16'h5555;
    LUT4 i26740_1_lut (.A(b[7]), .Z(n31879)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26740_1_lut.init = 16'h5555;
    LUT4 i26739_1_lut (.A(b[6]), .Z(n31878)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26739_1_lut.init = 16'h5555;
    LUT4 i26746_1_lut (.A(b[20]), .Z(n31885)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26746_1_lut.init = 16'h5555;
    LUT4 i26745_1_lut (.A(b[3]), .Z(n31884)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26745_1_lut.init = 16'h5555;
    LUT4 i26744_1_lut (.A(b[15]), .Z(n31883)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26744_1_lut.init = 16'h5555;
    LUT4 i26743_1_lut (.A(b[29]), .Z(n31882)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26743_1_lut.init = 16'h5555;
    LUT4 i26734_1_lut (.A(b[26]), .Z(n31873)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26734_1_lut.init = 16'h5555;
    LUT4 i26733_1_lut (.A(b[16]), .Z(n31872)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26733_1_lut.init = 16'h5555;
    LUT4 i26732_1_lut (.A(b[2]), .Z(n31871)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26732_1_lut.init = 16'h5555;
    LUT4 i26731_1_lut (.A(b[21]), .Z(n31870)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26731_1_lut.init = 16'h5555;
    LUT4 i26738_1_lut (.A(b[22]), .Z(n31877)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26738_1_lut.init = 16'h5555;
    LUT4 i26737_1_lut (.A(b[4]), .Z(n31876)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26737_1_lut.init = 16'h5555;
    LUT4 i26736_1_lut (.A(b[24]), .Z(n31875)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26736_1_lut.init = 16'h5555;
    LUT4 i26735_1_lut (.A(b[12]), .Z(n31874)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26735_1_lut.init = 16'h5555;
    LUT4 i26726_1_lut (.A(b[18]), .Z(n31865)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26726_1_lut.init = 16'h5555;
    LUT4 i26725_1_lut (.A(b[19]), .Z(n31864)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26725_1_lut.init = 16'h5555;
    LUT4 i26724_1_lut (.A(b[17]), .Z(n31863)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26724_1_lut.init = 16'h5555;
    LUT4 i26723_1_lut (.A(b[8]), .Z(n31862)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26723_1_lut.init = 16'h5555;
    LUT4 i26730_1_lut (.A(b[5]), .Z(n31869)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26730_1_lut.init = 16'h5555;
    LUT4 i26729_1_lut (.A(b[1]), .Z(n31868)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26729_1_lut.init = 16'h5555;
    LUT4 i26728_1_lut (.A(b[9]), .Z(n31867)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26728_1_lut.init = 16'h5555;
    LUT4 i26727_1_lut (.A(b[11]), .Z(n31866)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26727_1_lut.init = 16'h5555;
    LUT4 i26719_1_lut (.A(b[0]), .Z(n31858)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26719_1_lut.init = 16'h5555;
    LUT4 i26722_1_lut (.A(b[10]), .Z(n31861)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26722_1_lut.init = 16'h5555;
    LUT4 i26721_1_lut (.A(b[25]), .Z(n31860)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26721_1_lut.init = 16'h5555;
    LUT4 i26720_1_lut (.A(b[27]), .Z(n31859)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam i26720_1_lut.init = 16'h5555;
    LUT4 select_1205_Select_4_i1_3_lut_4_lut (.A(cycles[3]), .B(n41378), 
         .C(n41396), .D(cycles[4]), .Z(n1_adj_6191)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B !((D)+!C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(250[26:39])
    defparam select_1205_Select_4_i1_3_lut_4_lut.init = 16'he010;
    LUT4 i3333_2_lut_rep_1040 (.A(cycles[1]), .B(cycles[0]), .Z(n41445)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(250[26:39])
    defparam i3333_2_lut_rep_1040.init = 16'heeee;
    LUT4 i3341_2_lut_rep_973_3_lut (.A(cycles[1]), .B(cycles[0]), .C(cycles[2]), 
         .Z(n41378)) /* synthesis lut_function=(A+(B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(250[26:39])
    defparam i3341_2_lut_rep_973_3_lut.init = 16'hfefe;
    LUT4 i3349_2_lut_rep_888_3_lut_4_lut (.A(cycles[1]), .B(cycles[0]), 
         .C(cycles[3]), .D(cycles[2]), .Z(n41293)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(250[26:39])
    defparam i3349_2_lut_rep_888_3_lut_4_lut.init = 16'hfffe;
    LUT4 i4061_4_lut (.A(state[0]), .B(n32614), .C(divide_by_zero_x_N_3090), 
         .D(n15), .Z(n9351)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A ((D)+!B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i4061_4_lut.init = 16'h0ace;
    LUT4 i1_4_lut_adj_582 (.A(n41216), .B(n41196), .C(q_d), .D(n32608), 
         .Z(n32614)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_4_lut_adj_582.init = 16'h2000;
    LUT4 i4063_4_lut (.A(cycles_5__N_2934), .B(n9312), .C(n32658), .D(n15), 
         .Z(n9353)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i4063_4_lut.init = 16'heeec;
    LUT4 i1_4_lut_adj_583 (.A(n41196), .B(n41197), .C(n20863), .D(n32652), 
         .Z(n32658)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_583.init = 16'hfffe;
    
endmodule
//
// Verilog Description of module lm32_logic_op
//

module lm32_logic_op (\condition_x[2] , direction_x, operand_0_x, mc_result_x, 
            x_result_sel_mc_arith_x, logic_result_x, size_x, n36175, 
            n36178, n36184, n36190, n36193, n36196, n36199, n36223, 
            n36226, n36229, n36232, n36235, n36238, n36241, n36244, 
            n36247, n36250, n36253, n36256, n36259, n36262, n36265, 
            n36268, n36283, n36187) /* synthesis syn_module_defined=1 */ ;
    input \condition_x[2] ;
    input direction_x;
    input [31:0]operand_0_x;
    input [31:0]mc_result_x;
    input x_result_sel_mc_arith_x;
    output [31:0]logic_result_x;
    input [1:0]size_x;
    output n36175;
    output n36178;
    output n36184;
    output n36190;
    output n36193;
    output n36196;
    output n36199;
    output n36223;
    output n36226;
    output n36229;
    output n36232;
    output n36235;
    output n36238;
    output n36241;
    output n36244;
    output n36247;
    output n36250;
    output n36253;
    output n36256;
    output n36259;
    output n36262;
    output n36265;
    output n36268;
    output n36283;
    output n36187;
    
    
    wire n36188, n36284, n36269, n36266, n36263, n36260, n36257, 
        n36254, n36251, n36248, n36245, n36242, n36239, n36236, 
        n36233, n36230, n36227, n36224, n36200, n36197, n36194, 
        n36191, n36185, n36179, n36176, n36221, n36218, n36215, 
        n36212, n36209, n36206, n36203;
    
    LUT4 i31016_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[3]), 
         .Z(n36188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31016_3_lut.init = 16'hcaca;
    LUT4 i31112_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[31]), 
         .Z(n36284)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31112_3_lut.init = 16'hcaca;
    LUT4 i31097_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[30]), 
         .Z(n36269)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31097_3_lut.init = 16'hcaca;
    LUT4 i31094_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[29]), 
         .Z(n36266)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31094_3_lut.init = 16'hcaca;
    LUT4 i31091_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[28]), 
         .Z(n36263)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31091_3_lut.init = 16'hcaca;
    LUT4 i31088_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[27]), 
         .Z(n36260)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31088_3_lut.init = 16'hcaca;
    LUT4 i31085_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[26]), 
         .Z(n36257)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31085_3_lut.init = 16'hcaca;
    LUT4 i31082_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[25]), 
         .Z(n36254)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31082_3_lut.init = 16'hcaca;
    LUT4 i31079_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[24]), 
         .Z(n36251)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31079_3_lut.init = 16'hcaca;
    LUT4 i31076_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[23]), 
         .Z(n36248)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31076_3_lut.init = 16'hcaca;
    LUT4 i31073_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[22]), 
         .Z(n36245)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31073_3_lut.init = 16'hcaca;
    LUT4 i31070_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[21]), 
         .Z(n36242)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31070_3_lut.init = 16'hcaca;
    LUT4 i31067_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[20]), 
         .Z(n36239)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31067_3_lut.init = 16'hcaca;
    LUT4 i31064_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[19]), 
         .Z(n36236)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31064_3_lut.init = 16'hcaca;
    LUT4 i31061_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[18]), 
         .Z(n36233)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31061_3_lut.init = 16'hcaca;
    LUT4 i31058_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[17]), 
         .Z(n36230)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31058_3_lut.init = 16'hcaca;
    LUT4 i31055_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[16]), 
         .Z(n36227)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31055_3_lut.init = 16'hcaca;
    LUT4 i31052_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[15]), 
         .Z(n36224)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31052_3_lut.init = 16'hcaca;
    LUT4 i31028_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[7]), 
         .Z(n36200)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31028_3_lut.init = 16'hcaca;
    LUT4 i31025_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[6]), 
         .Z(n36197)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31025_3_lut.init = 16'hcaca;
    LUT4 i31022_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[5]), 
         .Z(n36194)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31022_3_lut.init = 16'hcaca;
    LUT4 i31019_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[4]), 
         .Z(n36191)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31019_3_lut.init = 16'hcaca;
    LUT4 i31013_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[2]), 
         .Z(n36185)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31013_3_lut.init = 16'hcaca;
    LUT4 i31007_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[1]), 
         .Z(n36179)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31007_3_lut.init = 16'hcaca;
    LUT4 i31004_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[0]), 
         .Z(n36176)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31004_3_lut.init = 16'hcaca;
    LUT4 i31050_3_lut (.A(n36221), .B(mc_result_x[14]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31050_3_lut.init = 16'hcaca;
    LUT4 i31049_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[14]), 
         .Z(n36221)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31049_3_lut.init = 16'hcaca;
    LUT4 i31047_3_lut (.A(n36218), .B(mc_result_x[13]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31047_3_lut.init = 16'hcaca;
    LUT4 i31046_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[13]), 
         .Z(n36218)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31046_3_lut.init = 16'hcaca;
    LUT4 i31044_3_lut (.A(n36215), .B(mc_result_x[12]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31044_3_lut.init = 16'hcaca;
    LUT4 i31043_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[12]), 
         .Z(n36215)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31043_3_lut.init = 16'hcaca;
    LUT4 i31041_3_lut (.A(n36212), .B(mc_result_x[11]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31041_3_lut.init = 16'hcaca;
    LUT4 i31040_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[11]), 
         .Z(n36212)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31040_3_lut.init = 16'hcaca;
    LUT4 i31038_3_lut (.A(n36209), .B(mc_result_x[10]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31038_3_lut.init = 16'hcaca;
    LUT4 i31037_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[10]), 
         .Z(n36209)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31037_3_lut.init = 16'hcaca;
    LUT4 i31035_3_lut (.A(n36206), .B(mc_result_x[9]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31035_3_lut.init = 16'hcaca;
    LUT4 i31034_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[9]), 
         .Z(n36206)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31034_3_lut.init = 16'hcaca;
    LUT4 i31032_3_lut (.A(n36203), .B(mc_result_x[8]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31032_3_lut.init = 16'hcaca;
    LUT4 i31031_3_lut (.A(\condition_x[2] ), .B(direction_x), .C(operand_0_x[8]), 
         .Z(n36203)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31031_3_lut.init = 16'hcaca;
    LUT4 i31003_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[0]), 
         .Z(n36175)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31003_3_lut.init = 16'hcaca;
    LUT4 i31006_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[1]), 
         .Z(n36178)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31006_3_lut.init = 16'hcaca;
    LUT4 i31012_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[2]), 
         .Z(n36184)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31012_3_lut.init = 16'hcaca;
    LUT4 i31018_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[4]), 
         .Z(n36190)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31018_3_lut.init = 16'hcaca;
    LUT4 i31021_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[5]), 
         .Z(n36193)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31021_3_lut.init = 16'hcaca;
    LUT4 i31024_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[6]), 
         .Z(n36196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31024_3_lut.init = 16'hcaca;
    LUT4 i31027_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[7]), 
         .Z(n36199)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31027_3_lut.init = 16'hcaca;
    LUT4 i31051_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[15]), 
         .Z(n36223)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31051_3_lut.init = 16'hcaca;
    LUT4 i31054_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[16]), 
         .Z(n36226)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31054_3_lut.init = 16'hcaca;
    LUT4 i31057_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[17]), 
         .Z(n36229)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31057_3_lut.init = 16'hcaca;
    LUT4 i31060_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[18]), 
         .Z(n36232)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31060_3_lut.init = 16'hcaca;
    LUT4 i31063_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[19]), 
         .Z(n36235)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31063_3_lut.init = 16'hcaca;
    LUT4 i31066_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[20]), 
         .Z(n36238)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31066_3_lut.init = 16'hcaca;
    LUT4 i31069_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[21]), 
         .Z(n36241)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31069_3_lut.init = 16'hcaca;
    LUT4 i31072_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[22]), 
         .Z(n36244)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31072_3_lut.init = 16'hcaca;
    LUT4 i31075_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[23]), 
         .Z(n36247)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31075_3_lut.init = 16'hcaca;
    LUT4 i31078_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[24]), 
         .Z(n36250)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31078_3_lut.init = 16'hcaca;
    LUT4 i31081_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[25]), 
         .Z(n36253)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31081_3_lut.init = 16'hcaca;
    LUT4 i31084_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[26]), 
         .Z(n36256)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31084_3_lut.init = 16'hcaca;
    LUT4 i31087_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[27]), 
         .Z(n36259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31087_3_lut.init = 16'hcaca;
    LUT4 i31090_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[28]), 
         .Z(n36262)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31090_3_lut.init = 16'hcaca;
    LUT4 i31093_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[29]), 
         .Z(n36265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31093_3_lut.init = 16'hcaca;
    LUT4 i31096_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[30]), 
         .Z(n36268)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31096_3_lut.init = 16'hcaca;
    LUT4 i31111_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[31]), 
         .Z(n36283)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31111_3_lut.init = 16'hcaca;
    LUT4 i31015_3_lut (.A(size_x[0]), .B(size_x[1]), .C(operand_0_x[3]), 
         .Z(n36187)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31015_3_lut.init = 16'hcaca;
    LUT4 i31005_3_lut (.A(n36176), .B(mc_result_x[0]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31005_3_lut.init = 16'hcaca;
    LUT4 i31008_3_lut (.A(n36179), .B(mc_result_x[1]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31008_3_lut.init = 16'hcaca;
    LUT4 i31014_3_lut (.A(n36185), .B(mc_result_x[2]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31014_3_lut.init = 16'hcaca;
    LUT4 i31020_3_lut (.A(n36191), .B(mc_result_x[4]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31020_3_lut.init = 16'hcaca;
    LUT4 i31023_3_lut (.A(n36194), .B(mc_result_x[5]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31023_3_lut.init = 16'hcaca;
    LUT4 i31026_3_lut (.A(n36197), .B(mc_result_x[6]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31026_3_lut.init = 16'hcaca;
    LUT4 i31029_3_lut (.A(n36200), .B(mc_result_x[7]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31029_3_lut.init = 16'hcaca;
    LUT4 i31053_3_lut (.A(n36224), .B(mc_result_x[15]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31053_3_lut.init = 16'hcaca;
    LUT4 i31056_3_lut (.A(n36227), .B(mc_result_x[16]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31056_3_lut.init = 16'hcaca;
    LUT4 i31059_3_lut (.A(n36230), .B(mc_result_x[17]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31059_3_lut.init = 16'hcaca;
    LUT4 i31062_3_lut (.A(n36233), .B(mc_result_x[18]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31062_3_lut.init = 16'hcaca;
    LUT4 i31065_3_lut (.A(n36236), .B(mc_result_x[19]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31065_3_lut.init = 16'hcaca;
    LUT4 i31068_3_lut (.A(n36239), .B(mc_result_x[20]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31068_3_lut.init = 16'hcaca;
    LUT4 i31071_3_lut (.A(n36242), .B(mc_result_x[21]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31071_3_lut.init = 16'hcaca;
    LUT4 i31074_3_lut (.A(n36245), .B(mc_result_x[22]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31074_3_lut.init = 16'hcaca;
    LUT4 i31077_3_lut (.A(n36248), .B(mc_result_x[23]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31077_3_lut.init = 16'hcaca;
    LUT4 i31080_3_lut (.A(n36251), .B(mc_result_x[24]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31080_3_lut.init = 16'hcaca;
    LUT4 i31083_3_lut (.A(n36254), .B(mc_result_x[25]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31083_3_lut.init = 16'hcaca;
    LUT4 i31086_3_lut (.A(n36257), .B(mc_result_x[26]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31086_3_lut.init = 16'hcaca;
    LUT4 i31089_3_lut (.A(n36260), .B(mc_result_x[27]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31089_3_lut.init = 16'hcaca;
    LUT4 i31092_3_lut (.A(n36263), .B(mc_result_x[28]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31092_3_lut.init = 16'hcaca;
    LUT4 i31095_3_lut (.A(n36266), .B(mc_result_x[29]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31095_3_lut.init = 16'hcaca;
    LUT4 i31098_3_lut (.A(n36269), .B(mc_result_x[30]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31098_3_lut.init = 16'hcaca;
    LUT4 i31113_3_lut (.A(n36284), .B(mc_result_x[31]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31113_3_lut.init = 16'hcaca;
    LUT4 i31017_3_lut (.A(n36188), .B(mc_result_x[3]), .C(x_result_sel_mc_arith_x), 
         .Z(logic_result_x[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i31017_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module \lm32_load_store_unit(base_address=32'b0,limit=32'b01111111111111111) 
//

module \lm32_load_store_unit(base_address=32'b0,limit=32'b01111111111111111)  (n41402, 
            \adder_result_x[1] , \adder_result_x[0] , n45171, n41283, 
            dcache_refill_request, n41215, REF_CLK_c, REF_CLK_c_enable_1235, 
            REF_CLK_c_enable_1606, size_x, LM32D_DAT_O, REF_CLK_c_enable_949, 
            REF_CLK_c_enable_1221, SHAREDBUS_DAT_O, LM32D_SEL_O, \LM32D_ADR_O[0] , 
            size_w, \LM32D_CTI_O[0] , n38965, \data_w[31] , \data_w[15] , 
            \operand_w[1] , stall_wb_load, \data_w[30] , \data_w[29] , 
            n30879, \data_w[28] , \data_w[27] , \data_w[26] , \data_w[25] , 
            \data_w[24] , store_operand_x, dcache_select_m, dcache_select_x, 
            wb_select_m, LM32D_STB_O, n41388, \condition_x[2] , LM32D_CYC_O, 
            REF_CLK_c_enable_1050, \load_data_w[16] , \load_data_w[17] , 
            \load_data_w[18] , \load_data_w[19] , \load_data_w[20] , \load_data_w[21] , 
            \load_data_w[22] , \load_data_w[23] , \load_data_w[24] , \load_data_w[25] , 
            \load_data_w[26] , \load_data_w[27] , \load_data_w[28] , \load_data_w[29] , 
            \load_data_w[30] , \load_data_w[31] , LM32D_WE_O, REF_CLK_c_enable_1234, 
            n12404, wb_load_complete, REF_CLK_c_enable_1236, n12400, 
            n21, \LM32D_ADR_O[1] , \LM32D_ADR_O[2] , \next_cycle_type[2] , 
            \LM32D_ADR_O[4] , \LM32D_ADR_O[5] , \d_adr_o_31__N_2278[5] , 
            \LM32D_ADR_O[6] , \LM32D_ADR_O[7] , \LM32D_ADR_O[8] , \LM32D_ADR_O[9] , 
            \d_adr_o_31__N_2278[9] , \LM32D_ADR_O[10] , \d_adr_o_31__N_2278[10] , 
            \LM32D_ADR_O[11] , \LM32D_ADR_O[12] , \LM32D_ADR_O[13] , \LM32D_ADR_O[14] , 
            \LM32D_ADR_O[15] , \LM32D_ADR_O[16] , \LM32D_ADR_O[17] , \LM32D_ADR_O[18] , 
            \LM32D_ADR_O[19] , \LM32D_ADR_O[20] , \LM32D_ADR_O[21] , \LM32D_ADR_O[22] , 
            \LM32D_ADR_O[23] , \LM32D_ADR_O[24] , \LM32D_ADR_O[25] , \d_adr_o_31__N_2278[25] , 
            \LM32D_ADR_O[26] , \LM32D_ADR_O[27] , \d_adr_o_31__N_2278[27] , 
            \LM32D_ADR_O[28] , \LM32D_ADR_O[29] , \LM32D_ADR_O[30] , \LM32D_ADR_O[31] , 
            REF_CLK_c_enable_1299, REF_CLK_c_enable_1304, \data_w[8] , 
            \data_w[9] , \data_w[10] , \data_w[11] , \data_w[12] , \data_w[13] , 
            \data_w[14] , \operand_w[0] , dcache_refilling, n41387, 
            n20639, n41380, locked_N_493, operand_m, n41217, exception_m, 
            n41232, n30070, n35745, n41233, n9, \load_data_w[6] , 
            n41144, n41145, n41156, n41157, n41140, n41141, n41164, 
            n41165, n41160, n41161, \load_data_w[7] , \load_data_w[5] , 
            \load_data_w[4] , n41148, n41149, \load_data_w[3] , n41152, 
            n41153, \load_data_w[2] , n41136, n41137, \load_data_w[1] , 
            \load_data_w[0] , icache_refill_request, n41435, branch_taken_m, 
            n41203, valid_d, q_d, n32652, \d_adr_o_31__N_2278[3] , 
            \d_adr_o_31__N_2278[2] , dcache_restart_request, n45183, state, 
            flush_set, flush_set_8__N_2513, \dcache_refill_address[5] , 
            \dcache_refill_address[9] , \dcache_refill_address[10] , \dcache_refill_address[25] , 
            \dcache_refill_address[27] , n41284, icache_restart_request, 
            n19852, valid_a, n30107, n9304, \state[2]_adj_192 , n41187, 
            n41196, n31996, n45175, way_match_0__N_2007, valid_f, 
            dflush_m, n41178, n36389, n37914, n37915, n37919, n37917, 
            n37916, n37918, n41, restart_request_N_1998, n15, n41172, 
            n32278, \tmem_write_address[1] , \tmem_write_address[5] , 
            \tmem_write_address[6] , n7502, VCC_net, GND_net, \genblk1.ra , 
            \dmem_write_address[3] , \dmem_write_address[7] , \dmem_write_address[8] , 
            n7388, n7322, n7256, n7204, n7190, n7206, n7208, \genblk1.ra_adj_202 , 
            n7224, n7222, n7220, n7356, n7354, n7352, n7350, n7348, 
            n7346, n7344, n7342, n7340, n7338, n7336, n7218, n7290, 
            n7288, n7286, n7284, n7216, n7282, n7280, n7278, n7214, 
            n7276, n7274, n7272, n7212, n7270, n7210) /* synthesis syn_module_defined=1 */ ;
    input n41402;
    input \adder_result_x[1] ;
    input \adder_result_x[0] ;
    input n45171;
    input n41283;
    output dcache_refill_request;
    input n41215;
    input REF_CLK_c;
    input REF_CLK_c_enable_1235;
    input REF_CLK_c_enable_1606;
    input [1:0]size_x;
    output [31:0]LM32D_DAT_O;
    input REF_CLK_c_enable_949;
    input REF_CLK_c_enable_1221;
    input [31:0]SHAREDBUS_DAT_O;
    output [3:0]LM32D_SEL_O;
    output \LM32D_ADR_O[0] ;
    output [1:0]size_w;
    output \LM32D_CTI_O[0] ;
    input n38965;
    output \data_w[31] ;
    output \data_w[15] ;
    input \operand_w[1] ;
    output stall_wb_load;
    output \data_w[30] ;
    output \data_w[29] ;
    input n30879;
    output \data_w[28] ;
    output \data_w[27] ;
    output \data_w[26] ;
    output \data_w[25] ;
    output \data_w[24] ;
    input [31:0]store_operand_x;
    output dcache_select_m;
    input dcache_select_x;
    output wb_select_m;
    output LM32D_STB_O;
    input n41388;
    input \condition_x[2] ;
    output LM32D_CYC_O;
    input REF_CLK_c_enable_1050;
    output \load_data_w[16] ;
    output \load_data_w[17] ;
    output \load_data_w[18] ;
    output \load_data_w[19] ;
    output \load_data_w[20] ;
    output \load_data_w[21] ;
    output \load_data_w[22] ;
    output \load_data_w[23] ;
    output \load_data_w[24] ;
    output \load_data_w[25] ;
    output \load_data_w[26] ;
    output \load_data_w[27] ;
    output \load_data_w[28] ;
    output \load_data_w[29] ;
    output \load_data_w[30] ;
    output \load_data_w[31] ;
    output LM32D_WE_O;
    input REF_CLK_c_enable_1234;
    input n12404;
    output wb_load_complete;
    input REF_CLK_c_enable_1236;
    input n12400;
    output n21;
    output \LM32D_ADR_O[1] ;
    output \LM32D_ADR_O[2] ;
    output \next_cycle_type[2] ;
    output \LM32D_ADR_O[4] ;
    output \LM32D_ADR_O[5] ;
    input \d_adr_o_31__N_2278[5] ;
    output \LM32D_ADR_O[6] ;
    output \LM32D_ADR_O[7] ;
    output \LM32D_ADR_O[8] ;
    output \LM32D_ADR_O[9] ;
    input \d_adr_o_31__N_2278[9] ;
    output \LM32D_ADR_O[10] ;
    input \d_adr_o_31__N_2278[10] ;
    output \LM32D_ADR_O[11] ;
    output \LM32D_ADR_O[12] ;
    output \LM32D_ADR_O[13] ;
    output \LM32D_ADR_O[14] ;
    output \LM32D_ADR_O[15] ;
    output \LM32D_ADR_O[16] ;
    output \LM32D_ADR_O[17] ;
    output \LM32D_ADR_O[18] ;
    output \LM32D_ADR_O[19] ;
    output \LM32D_ADR_O[20] ;
    output \LM32D_ADR_O[21] ;
    output \LM32D_ADR_O[22] ;
    output \LM32D_ADR_O[23] ;
    output \LM32D_ADR_O[24] ;
    output \LM32D_ADR_O[25] ;
    input \d_adr_o_31__N_2278[25] ;
    output \LM32D_ADR_O[26] ;
    output \LM32D_ADR_O[27] ;
    input \d_adr_o_31__N_2278[27] ;
    output \LM32D_ADR_O[28] ;
    output \LM32D_ADR_O[29] ;
    output \LM32D_ADR_O[30] ;
    output \LM32D_ADR_O[31] ;
    input REF_CLK_c_enable_1299;
    input REF_CLK_c_enable_1304;
    output \data_w[8] ;
    output \data_w[9] ;
    output \data_w[10] ;
    output \data_w[11] ;
    output \data_w[12] ;
    output \data_w[13] ;
    output \data_w[14] ;
    input \operand_w[0] ;
    output dcache_refilling;
    output n41387;
    output n20639;
    input n41380;
    input locked_N_493;
    input [31:0]operand_m;
    input n41217;
    input exception_m;
    input n41232;
    input n30070;
    input n35745;
    input n41233;
    input n9;
    output \load_data_w[6] ;
    input n41144;
    output n41145;
    input n41156;
    output n41157;
    input n41140;
    output n41141;
    input n41164;
    output n41165;
    input n41160;
    output n41161;
    output \load_data_w[7] ;
    output \load_data_w[5] ;
    output \load_data_w[4] ;
    input n41148;
    output n41149;
    output \load_data_w[3] ;
    input n41152;
    output n41153;
    output \load_data_w[2] ;
    input n41136;
    output n41137;
    output \load_data_w[1] ;
    output \load_data_w[0] ;
    input icache_refill_request;
    output n41435;
    input branch_taken_m;
    output n41203;
    input valid_d;
    output q_d;
    output n32652;
    input \d_adr_o_31__N_2278[3] ;
    input \d_adr_o_31__N_2278[2] ;
    output dcache_restart_request;
    input n45183;
    output [2:0]state;
    output [8:0]flush_set;
    input [8:0]flush_set_8__N_2513;
    output \dcache_refill_address[5] ;
    output \dcache_refill_address[9] ;
    output \dcache_refill_address[10] ;
    output \dcache_refill_address[25] ;
    output \dcache_refill_address[27] ;
    input n41284;
    input icache_restart_request;
    input n19852;
    output valid_a;
    input n30107;
    input n9304;
    input \state[2]_adj_192 ;
    input n41187;
    input n41196;
    output n31996;
    input n45175;
    input way_match_0__N_2007;
    input valid_f;
    input dflush_m;
    output n41178;
    output n36389;
    output n37914;
    output n37915;
    output n37919;
    output n37917;
    output n37916;
    output n37918;
    input n41;
    output restart_request_N_1998;
    input n15;
    output n41172;
    output n32278;
    input \tmem_write_address[1] ;
    input \tmem_write_address[5] ;
    input \tmem_write_address[6] ;
    input [8:0]n7502;
    input VCC_net;
    input GND_net;
    output [8:0]\genblk1.ra ;
    input \dmem_write_address[3] ;
    input \dmem_write_address[7] ;
    input \dmem_write_address[8] ;
    input [10:0]n7388;
    input [10:0]n7322;
    input [10:0]n7256;
    output n7204;
    input [10:0]n7190;
    output n7206;
    output n7208;
    output [10:0]\genblk1.ra_adj_202 ;
    output n7224;
    output n7222;
    output n7220;
    output n7356;
    output n7354;
    output n7352;
    output n7350;
    output n7348;
    output n7346;
    output n7344;
    output n7342;
    output n7340;
    output n7338;
    output n7336;
    output n7218;
    output n7290;
    output n7288;
    output n7286;
    output n7284;
    output n7216;
    output n7282;
    output n7280;
    output n7278;
    output n7214;
    output n7276;
    output n7274;
    output n7272;
    output n7212;
    output n7270;
    output n7210;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    
    wire n9_c;
    wire [3:0]byte_enable_x;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(245[29:42])
    
    wire n11;
    wire [1:0]size_m;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(239[22:28])
    wire [31:0]store_data_m;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(244[22:34])
    wire [31:0]wb_data_m;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(276[22:31])
    
    wire REF_CLK_c_enable_1270;
    wire [3:0]d_sel_o_3__N_2358;
    wire [31:0]d_adr_o_31__N_2278;
    wire [3:0]byte_enable_m;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(246[29:42])
    wire [31:0]store_data_x;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(243[22:34])
    wire [31:0]data_w;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(248[22:28])
    wire [31:0]data_m;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(247[23:29])
    
    wire REF_CLK_c_enable_1242, sign_extend_w, sign_extend_m, n35;
    wire [1:0]size_w_c;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(240[22:28])
    
    wire n32, n34758, n27, REF_CLK_c_enable_193, n31463, n32_adj_6042, 
        n32_adj_6043, dcache_refill_ready, n32_adj_6044, n32_adj_6045, 
        n32_adj_6046, n32_adj_6047, n32_adj_6048, n32_adj_6049, n32_adj_6050, 
        n32_adj_6051, n32_adj_6052, n32_adj_6053, n32_adj_6054, n32_adj_6055, 
        n32_adj_6056, dcache_select_x_N_2440, REF_CLK_c_enable_398, n12384, 
        n23, n28, n31, n23_adj_6057, n28_adj_6058, n31_adj_6059, 
        n23_adj_6060, n28_adj_6061, n31_adj_6062, n23_adj_6063, n28_adj_6064, 
        n31_adj_6065, n23_adj_6066, n28_adj_6067, n31_adj_6068, n23_adj_6069, 
        n28_adj_6070, n31_adj_6071, n20800, n41489, n41490, n23_adj_6072, 
        n28_adj_6073, n31_adj_6074, n23_adj_6075, n28_adj_6076, n31_adj_6077, 
        n25, n25_adj_6078, n25_adj_6079, n25_adj_6080, n25_adj_6081, 
        n25_adj_6082, n25_adj_6083;
    wire [31:0]d_adr_o_31__N_2149;
    
    wire n32298;
    wire [1:0]n3722;
    wire [31:0]dcache_refill_address;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(254[23:44])
    
    wire n2, n2_adj_6084, n2_adj_6085, n2_adj_6086, n2_adj_6087, n2_adj_6088, 
        n2_adj_6089, n2_adj_6090;
    wire [7:0]dcache_data_m;
    wire [7:0]n6416;
    wire [7:0]n6417;
    
    wire n41392, n35694;
    wire [7:0]n6418;
    
    wire n34978, n25_adj_6092;
    
    LUT4 i1_3_lut_4_lut (.A(n41402), .B(\adder_result_x[1] ), .C(n9_c), 
         .D(\adder_result_x[0] ), .Z(byte_enable_x[0])) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(461[5:29])
    defparam i1_3_lut_4_lut.init = 16'hf4f0;
    LUT4 i1_3_lut_4_lut_adj_436 (.A(n41402), .B(\adder_result_x[1] ), .C(n9_c), 
         .D(\adder_result_x[0] ), .Z(byte_enable_x[1])) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(461[5:29])
    defparam i1_3_lut_4_lut_adj_436.init = 16'hf0f4;
    LUT4 i1_3_lut_4_lut_adj_437 (.A(n45171), .B(n41283), .C(dcache_refill_request), 
         .D(n41215), .Z(n11)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i1_3_lut_4_lut_adj_437.init = 16'hfff8;
    FD1P3DX size_m_i0_i0 (.D(size_x[0]), .SP(REF_CLK_c_enable_1235), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(size_m[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam size_m_i0_i0.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i0 (.D(store_data_m[0]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i0.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i0 (.D(SHAREDBUS_DAT_O[0]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i0.GSR = "ENABLED";
    FD1P3DX d_sel_o_i0_i0 (.D(d_sel_o_3__N_2358[0]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_SEL_O[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_sel_o_i0_i0.GSR = "ENABLED";
    FD1P3DX d_adr_o_i0 (.D(d_adr_o_31__N_2278[0]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[0] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0.GSR = "ENABLED";
    FD1P3DX byte_enable_m_i0_i0 (.D(byte_enable_x[0]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(byte_enable_m[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam byte_enable_m_i0_i0.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i0 (.D(store_data_x[0]), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i0.GSR = "ENABLED";
    FD1S3DX size_w_i0 (.D(size_m[0]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(size_w[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam size_w_i0.GSR = "ENABLED";
    FD1S3DX data_w_i0 (.D(data_m[0]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(data_w[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i0.GSR = "ENABLED";
    FD1P3BX d_cti_o_i0 (.D(n38965), .SP(REF_CLK_c_enable_1242), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(\LM32D_CTI_O[0] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_cti_o_i0.GSR = "ENABLED";
    FD1S3DX sign_extend_w_183 (.D(sign_extend_m), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(sign_extend_w)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam sign_extend_w_183.GSR = "ENABLED";
    LUT4 i56_3_lut (.A(n35), .B(\data_w[31] ), .C(size_w_c[1]), .Z(n32)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(n34758), .B(\data_w[31] ), .C(\data_w[15] ), .D(\operand_w[1] ), 
         .Z(n27)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut.init = 16'ha088;
    LUT4 i1_2_lut (.A(size_w_c[1]), .B(sign_extend_w), .Z(n34758)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_2_lut.init = 16'h8888;
    FD1P3DX stall_wb_load_173 (.D(n31463), .SP(REF_CLK_c_enable_193), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(stall_wb_load)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam stall_wb_load_173.GSR = "ENABLED";
    LUT4 i56_3_lut_adj_438 (.A(n35), .B(\data_w[30] ), .C(size_w_c[1]), 
         .Z(n32_adj_6042)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_438.init = 16'hcaca;
    LUT4 i56_3_lut_adj_439 (.A(n35), .B(\data_w[29] ), .C(size_w_c[1]), 
         .Z(n32_adj_6043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_439.init = 16'hcaca;
    FD1S3DX dcache_refill_ready_174 (.D(n30879), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(dcache_refill_ready)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam dcache_refill_ready_174.GSR = "ENABLED";
    LUT4 i56_3_lut_adj_440 (.A(n35), .B(\data_w[28] ), .C(size_w_c[1]), 
         .Z(n32_adj_6044)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_440.init = 16'hcaca;
    LUT4 i56_3_lut_adj_441 (.A(n35), .B(\data_w[27] ), .C(size_w_c[1]), 
         .Z(n32_adj_6045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_441.init = 16'hcaca;
    LUT4 i56_3_lut_adj_442 (.A(n35), .B(\data_w[26] ), .C(size_w_c[1]), 
         .Z(n32_adj_6046)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_442.init = 16'hcaca;
    LUT4 i56_3_lut_adj_443 (.A(n35), .B(\data_w[25] ), .C(size_w_c[1]), 
         .Z(n32_adj_6047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_443.init = 16'hcaca;
    LUT4 i56_3_lut_adj_444 (.A(n35), .B(\data_w[24] ), .C(size_w_c[1]), 
         .Z(n32_adj_6048)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_444.init = 16'hcaca;
    LUT4 i56_3_lut_adj_445 (.A(n35), .B(data_w[23]), .C(size_w_c[1]), 
         .Z(n32_adj_6049)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_445.init = 16'hcaca;
    LUT4 i56_3_lut_adj_446 (.A(n35), .B(data_w[22]), .C(size_w_c[1]), 
         .Z(n32_adj_6050)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_446.init = 16'hcaca;
    LUT4 i56_3_lut_adj_447 (.A(n35), .B(data_w[21]), .C(size_w_c[1]), 
         .Z(n32_adj_6051)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_447.init = 16'hcaca;
    LUT4 i56_3_lut_adj_448 (.A(n35), .B(data_w[20]), .C(size_w_c[1]), 
         .Z(n32_adj_6052)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_448.init = 16'hcaca;
    LUT4 i56_3_lut_adj_449 (.A(n35), .B(data_w[19]), .C(size_w_c[1]), 
         .Z(n32_adj_6053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_449.init = 16'hcaca;
    LUT4 i56_3_lut_adj_450 (.A(n35), .B(data_w[18]), .C(size_w_c[1]), 
         .Z(n32_adj_6054)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_450.init = 16'hcaca;
    LUT4 i56_3_lut_adj_451 (.A(n35), .B(data_w[17]), .C(size_w_c[1]), 
         .Z(n32_adj_6055)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_451.init = 16'hcaca;
    LUT4 i56_3_lut_adj_452 (.A(n35), .B(data_w[16]), .C(size_w_c[1]), 
         .Z(n32_adj_6056)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_452.init = 16'hcaca;
    LUT4 store_operand_x_0__bdd_4_lut (.A(store_operand_x[0]), .B(size_x[1]), 
         .C(store_operand_x[16]), .D(size_x[0]), .Z(store_data_x[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(((D)+!C)+!B)) */ ;
    defparam store_operand_x_0__bdd_4_lut.init = 16'h88e2;
    LUT4 store_operand_x_1__bdd_4_lut (.A(store_operand_x[1]), .B(size_x[1]), 
         .C(store_operand_x[17]), .D(size_x[0]), .Z(store_data_x[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(((D)+!C)+!B)) */ ;
    defparam store_operand_x_1__bdd_4_lut.init = 16'h88e2;
    LUT4 store_operand_x_2__bdd_4_lut (.A(store_operand_x[2]), .B(size_x[1]), 
         .C(store_operand_x[18]), .D(size_x[0]), .Z(store_data_x[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(((D)+!C)+!B)) */ ;
    defparam store_operand_x_2__bdd_4_lut.init = 16'h88e2;
    LUT4 store_operand_x_3__bdd_4_lut (.A(store_operand_x[3]), .B(size_x[1]), 
         .C(store_operand_x[19]), .D(size_x[0]), .Z(store_data_x[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(((D)+!C)+!B)) */ ;
    defparam store_operand_x_3__bdd_4_lut.init = 16'h88e2;
    LUT4 store_operand_x_7__bdd_4_lut (.A(store_operand_x[7]), .B(size_x[1]), 
         .C(store_operand_x[23]), .D(size_x[0]), .Z(store_data_x[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(((D)+!C)+!B)) */ ;
    defparam store_operand_x_7__bdd_4_lut.init = 16'h88e2;
    LUT4 store_operand_x_6__bdd_4_lut (.A(store_operand_x[6]), .B(size_x[1]), 
         .C(store_operand_x[22]), .D(size_x[0]), .Z(store_data_x[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(((D)+!C)+!B)) */ ;
    defparam store_operand_x_6__bdd_4_lut.init = 16'h88e2;
    FD1P3DX dcache_select_m_179 (.D(dcache_select_x), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(dcache_select_m)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam dcache_select_m_179.GSR = "ENABLED";
    FD1P3DX wb_select_m_180 (.D(dcache_select_x_N_2440), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_select_m)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam wb_select_m_180.GSR = "ENABLED";
    FD1P3DX d_stb_o_163 (.D(n41388), .SP(REF_CLK_c_enable_398), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(LM32D_STB_O)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_stb_o_163.GSR = "ENABLED";
    LUT4 store_operand_x_4__bdd_4_lut (.A(store_operand_x[4]), .B(size_x[1]), 
         .C(store_operand_x[20]), .D(size_x[0]), .Z(store_data_x[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(((D)+!C)+!B)) */ ;
    defparam store_operand_x_4__bdd_4_lut.init = 16'h88e2;
    LUT4 store_operand_x_5__bdd_4_lut (.A(store_operand_x[5]), .B(size_x[1]), 
         .C(store_operand_x[21]), .D(size_x[0]), .Z(store_data_x[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(((D)+!C)+!B)) */ ;
    defparam store_operand_x_5__bdd_4_lut.init = 16'h88e2;
    FD1P3DX sign_extend_m_175 (.D(\condition_x[2] ), .SP(REF_CLK_c_enable_1235), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(sign_extend_m)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam sign_extend_m_175.GSR = "ENABLED";
    FD1S3DX d_cyc_o_162 (.D(n12384), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(LM32D_CYC_O)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_cyc_o_162.GSR = "ENABLED";
    PFUMX i52 (.BLUT(n23), .ALUT(n28), .C0(\operand_w[1] ), .Z(n31));
    PFUMX i52_adj_453 (.BLUT(n23_adj_6057), .ALUT(n28_adj_6058), .C0(\operand_w[1] ), 
          .Z(n31_adj_6059));
    PFUMX i52_adj_454 (.BLUT(n23_adj_6060), .ALUT(n28_adj_6061), .C0(\operand_w[1] ), 
          .Z(n31_adj_6062));
    PFUMX i52_adj_455 (.BLUT(n23_adj_6063), .ALUT(n28_adj_6064), .C0(\operand_w[1] ), 
          .Z(n31_adj_6065));
    PFUMX i52_adj_456 (.BLUT(n23_adj_6066), .ALUT(n28_adj_6067), .C0(\operand_w[1] ), 
          .Z(n31_adj_6068));
    PFUMX i52_adj_457 (.BLUT(n23_adj_6069), .ALUT(n28_adj_6070), .C0(\operand_w[1] ), 
          .Z(n31_adj_6071));
    LUT4 i1_3_lut_4_lut_adj_458 (.A(n41402), .B(\adder_result_x[1] ), .C(n20800), 
         .D(\adder_result_x[0] ), .Z(byte_enable_x[2])) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !((D)+!C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(463[5:29])
    defparam i1_3_lut_4_lut_adj_458.init = 16'h1f0f;
    FD1P3DX size_m_i0_i1 (.D(size_x[1]), .SP(REF_CLK_c_enable_1050), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(size_m[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam size_m_i0_i1.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i1 (.D(store_data_m[1]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i1.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i2 (.D(store_data_m[2]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i2.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i3 (.D(store_data_m[3]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i3.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i4 (.D(store_data_m[4]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i4.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i5 (.D(store_data_m[5]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i5.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i6 (.D(store_data_m[6]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i6.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i7 (.D(store_data_m[7]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i7.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i8 (.D(store_data_m[8]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i8.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i9 (.D(store_data_m[9]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i9.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i10 (.D(store_data_m[10]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i10.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i11 (.D(store_data_m[11]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i11.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i12 (.D(store_data_m[12]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i12.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i13 (.D(store_data_m[13]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i13.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i14 (.D(store_data_m[14]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i14.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i15 (.D(store_data_m[15]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i15.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i16 (.D(store_data_m[16]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i16.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i17 (.D(store_data_m[17]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i17.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i18 (.D(store_data_m[18]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i18.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i19 (.D(store_data_m[19]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i19.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i20 (.D(store_data_m[20]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i20.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i21 (.D(store_data_m[21]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i21.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i22 (.D(store_data_m[22]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i22.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i23 (.D(store_data_m[23]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i23.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i24 (.D(store_data_m[24]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i24.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i25 (.D(store_data_m[25]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i25.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i26 (.D(store_data_m[26]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i26.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i27 (.D(store_data_m[27]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i27.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i28 (.D(store_data_m[28]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i28.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i29 (.D(store_data_m[29]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i29.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i30 (.D(store_data_m[30]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i30.GSR = "ENABLED";
    FD1P3DX d_dat_o_i0_i31 (.D(store_data_m[31]), .SP(REF_CLK_c_enable_949), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_DAT_O[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i31.GSR = "ENABLED";
    LUT4 i33226_3_lut_4_lut (.A(n41402), .B(\adder_result_x[1] ), .C(n20800), 
         .D(\adder_result_x[0] ), .Z(byte_enable_x[3])) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(463[5:29])
    defparam i33226_3_lut_4_lut.init = 16'h0f1f;
    PFUMX i34379 (.BLUT(n41489), .ALUT(n41490), .C0(\operand_w[1] ), .Z(n35));
    PFUMX i52_adj_459 (.BLUT(n23_adj_6072), .ALUT(n28_adj_6073), .C0(\operand_w[1] ), 
          .Z(n31_adj_6074));
    PFUMX i52_adj_460 (.BLUT(n23_adj_6075), .ALUT(n28_adj_6076), .C0(\operand_w[1] ), 
          .Z(n31_adj_6077));
    LUT4 i55_3_lut (.A(n32_adj_6056), .B(n27), .C(size_w[0]), .Z(\load_data_w[16] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut.init = 16'hcaca;
    LUT4 i55_3_lut_adj_461 (.A(n32_adj_6055), .B(n27), .C(size_w[0]), 
         .Z(\load_data_w[17] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_461.init = 16'hcaca;
    LUT4 i55_3_lut_adj_462 (.A(n32_adj_6054), .B(n27), .C(size_w[0]), 
         .Z(\load_data_w[18] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_462.init = 16'hcaca;
    LUT4 i55_3_lut_adj_463 (.A(n32_adj_6053), .B(n27), .C(size_w[0]), 
         .Z(\load_data_w[19] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_463.init = 16'hcaca;
    LUT4 i55_3_lut_adj_464 (.A(n32_adj_6052), .B(n27), .C(size_w[0]), 
         .Z(\load_data_w[20] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_464.init = 16'hcaca;
    LUT4 i55_3_lut_adj_465 (.A(n32_adj_6051), .B(n27), .C(size_w[0]), 
         .Z(\load_data_w[21] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_465.init = 16'hcaca;
    FD1P3DX wb_data_m_i0_i1 (.D(SHAREDBUS_DAT_O[1]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i1.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i2 (.D(SHAREDBUS_DAT_O[2]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i2.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i3 (.D(SHAREDBUS_DAT_O[3]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i3.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i4 (.D(SHAREDBUS_DAT_O[4]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i4.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i5 (.D(SHAREDBUS_DAT_O[5]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i5.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i6 (.D(SHAREDBUS_DAT_O[6]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i6.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i7 (.D(SHAREDBUS_DAT_O[7]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i7.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i8 (.D(SHAREDBUS_DAT_O[8]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i8.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i9 (.D(SHAREDBUS_DAT_O[9]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i9.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i10 (.D(SHAREDBUS_DAT_O[10]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i10.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i11 (.D(SHAREDBUS_DAT_O[11]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i11.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i12 (.D(SHAREDBUS_DAT_O[12]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i12.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i13 (.D(SHAREDBUS_DAT_O[13]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i13.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i14 (.D(SHAREDBUS_DAT_O[14]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i14.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i15 (.D(SHAREDBUS_DAT_O[15]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i15.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i16 (.D(SHAREDBUS_DAT_O[16]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i16.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i17 (.D(SHAREDBUS_DAT_O[17]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i17.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i18 (.D(SHAREDBUS_DAT_O[18]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i18.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i19 (.D(SHAREDBUS_DAT_O[19]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i19.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i20 (.D(SHAREDBUS_DAT_O[20]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i20.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i21 (.D(SHAREDBUS_DAT_O[21]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i21.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i22 (.D(SHAREDBUS_DAT_O[22]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i22.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i23 (.D(SHAREDBUS_DAT_O[23]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i23.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i24 (.D(SHAREDBUS_DAT_O[24]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i24.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i25 (.D(SHAREDBUS_DAT_O[25]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i25.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i26 (.D(SHAREDBUS_DAT_O[26]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i26.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i27 (.D(SHAREDBUS_DAT_O[27]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i27.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i28 (.D(SHAREDBUS_DAT_O[28]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i28.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i29 (.D(SHAREDBUS_DAT_O[29]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i29.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i30 (.D(SHAREDBUS_DAT_O[30]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i30.GSR = "ENABLED";
    FD1P3DX wb_data_m_i0_i31 (.D(SHAREDBUS_DAT_O[31]), .SP(REF_CLK_c_enable_1221), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_data_m[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i31.GSR = "ENABLED";
    FD1P3DX d_sel_o_i0_i1 (.D(d_sel_o_3__N_2358[1]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_SEL_O[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_sel_o_i0_i1.GSR = "ENABLED";
    LUT4 i55_3_lut_adj_466 (.A(n32_adj_6050), .B(n27), .C(size_w[0]), 
         .Z(\load_data_w[22] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_466.init = 16'hcaca;
    LUT4 i55_3_lut_adj_467 (.A(n32_adj_6049), .B(n27), .C(size_w[0]), 
         .Z(\load_data_w[23] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_467.init = 16'hcaca;
    LUT4 i55_3_lut_adj_468 (.A(n32_adj_6048), .B(n27), .C(size_w[0]), 
         .Z(\load_data_w[24] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_468.init = 16'hcaca;
    LUT4 i55_3_lut_adj_469 (.A(n32_adj_6047), .B(n27), .C(size_w[0]), 
         .Z(\load_data_w[25] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_469.init = 16'hcaca;
    LUT4 i55_3_lut_adj_470 (.A(n32_adj_6046), .B(n27), .C(size_w[0]), 
         .Z(\load_data_w[26] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_470.init = 16'hcaca;
    LUT4 i55_3_lut_adj_471 (.A(n32_adj_6045), .B(n27), .C(size_w[0]), 
         .Z(\load_data_w[27] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_471.init = 16'hcaca;
    LUT4 i55_3_lut_adj_472 (.A(n32_adj_6044), .B(n27), .C(size_w[0]), 
         .Z(\load_data_w[28] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_472.init = 16'hcaca;
    LUT4 i55_3_lut_adj_473 (.A(n32_adj_6043), .B(n27), .C(size_w[0]), 
         .Z(\load_data_w[29] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_473.init = 16'hcaca;
    LUT4 i55_3_lut_adj_474 (.A(n32_adj_6042), .B(n27), .C(size_w[0]), 
         .Z(\load_data_w[30] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_474.init = 16'hcaca;
    LUT4 i55_3_lut_adj_475 (.A(n32), .B(n27), .C(size_w[0]), .Z(\load_data_w[31] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_475.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut (.A(data_w[17]), .B(data_w[1]), .C(\operand_w[1] ), 
         .D(size_w[0]), .Z(n25)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut.init = 16'hcacc;
    LUT4 i1_4_lut_4_lut_adj_476 (.A(data_w[18]), .B(data_w[2]), .C(\operand_w[1] ), 
         .D(size_w[0]), .Z(n25_adj_6078)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_476.init = 16'hcacc;
    LUT4 i1_4_lut_4_lut_adj_477 (.A(data_w[19]), .B(data_w[3]), .C(\operand_w[1] ), 
         .D(size_w[0]), .Z(n25_adj_6079)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_477.init = 16'hcacc;
    LUT4 i1_4_lut_4_lut_adj_478 (.A(data_w[20]), .B(data_w[4]), .C(\operand_w[1] ), 
         .D(size_w[0]), .Z(n25_adj_6080)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_478.init = 16'hcacc;
    FD1P3DX d_we_o_167 (.D(n12404), .SP(REF_CLK_c_enable_1234), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(LM32D_WE_O)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_we_o_167.GSR = "ENABLED";
    FD1P3DX wb_load_complete_172 (.D(n12400), .SP(REF_CLK_c_enable_1236), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(wb_load_complete)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_load_complete_172.GSR = "ENABLED";
    LUT4 i1_4_lut_4_lut_adj_479 (.A(data_w[21]), .B(data_w[5]), .C(\operand_w[1] ), 
         .D(size_w[0]), .Z(n25_adj_6081)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_479.init = 16'hcacc;
    LUT4 i1_4_lut_4_lut_adj_480 (.A(data_w[22]), .B(data_w[6]), .C(\operand_w[1] ), 
         .D(size_w[0]), .Z(n25_adj_6082)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_480.init = 16'hcacc;
    LUT4 i1_4_lut_4_lut_adj_481 (.A(data_w[23]), .B(data_w[7]), .C(\operand_w[1] ), 
         .D(size_w[0]), .Z(n25_adj_6083)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_481.init = 16'hcacc;
    LUT4 i1_2_lut_adj_482 (.A(LM32D_SEL_O[0]), .B(LM32D_SEL_O[1]), .Z(n21)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_482.init = 16'h8888;
    FD1P3DX d_sel_o_i0_i2 (.D(d_sel_o_3__N_2358[2]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_SEL_O[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_sel_o_i0_i2.GSR = "ENABLED";
    FD1P3DX d_sel_o_i0_i3 (.D(d_sel_o_3__N_2358[3]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(LM32D_SEL_O[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_sel_o_i0_i3.GSR = "ENABLED";
    FD1P3DX d_adr_o_i1 (.D(d_adr_o_31__N_2278[1]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[1] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i1.GSR = "ENABLED";
    FD1P3DX d_adr_o_i2 (.D(d_adr_o_31__N_2149[2]), .SP(REF_CLK_c_enable_1242), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i2.GSR = "ENABLED";
    FD1P3DX d_adr_o_i3 (.D(d_adr_o_31__N_2149[3]), .SP(REF_CLK_c_enable_1242), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\next_cycle_type[2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i3.GSR = "ENABLED";
    FD1P3DX d_adr_o_i4 (.D(d_adr_o_31__N_2278[4]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i4.GSR = "ENABLED";
    FD1P3DX d_adr_o_i5 (.D(\d_adr_o_31__N_2278[5] ), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[5] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i5.GSR = "ENABLED";
    FD1P3DX d_adr_o_i6 (.D(d_adr_o_31__N_2278[6]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[6] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i6.GSR = "ENABLED";
    FD1P3DX d_adr_o_i7 (.D(d_adr_o_31__N_2278[7]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[7] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i7.GSR = "ENABLED";
    FD1P3DX d_adr_o_i8 (.D(d_adr_o_31__N_2278[8]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[8] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i8.GSR = "ENABLED";
    FD1P3DX d_adr_o_i9 (.D(\d_adr_o_31__N_2278[9] ), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[9] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i9.GSR = "ENABLED";
    FD1P3DX d_adr_o_i10 (.D(\d_adr_o_31__N_2278[10] ), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[10] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i10.GSR = "ENABLED";
    FD1P3DX d_adr_o_i11 (.D(d_adr_o_31__N_2278[11]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[11] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i11.GSR = "ENABLED";
    FD1P3DX d_adr_o_i12 (.D(d_adr_o_31__N_2278[12]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[12] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i12.GSR = "ENABLED";
    FD1P3DX d_adr_o_i13 (.D(d_adr_o_31__N_2278[13]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[13] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i13.GSR = "ENABLED";
    FD1P3DX d_adr_o_i14 (.D(d_adr_o_31__N_2278[14]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[14] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i14.GSR = "ENABLED";
    FD1P3DX d_adr_o_i15 (.D(d_adr_o_31__N_2278[15]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[15] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i15.GSR = "ENABLED";
    FD1P3DX d_adr_o_i16 (.D(d_adr_o_31__N_2278[16]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[16] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i16.GSR = "ENABLED";
    FD1P3DX d_adr_o_i17 (.D(d_adr_o_31__N_2278[17]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[17] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i17.GSR = "ENABLED";
    FD1P3DX d_adr_o_i18 (.D(d_adr_o_31__N_2278[18]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[18] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i18.GSR = "ENABLED";
    FD1P3DX d_adr_o_i19 (.D(d_adr_o_31__N_2278[19]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[19] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i19.GSR = "ENABLED";
    FD1P3DX d_adr_o_i20 (.D(d_adr_o_31__N_2278[20]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[20] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i20.GSR = "ENABLED";
    FD1P3DX d_adr_o_i21 (.D(d_adr_o_31__N_2278[21]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[21] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i21.GSR = "ENABLED";
    FD1P3DX d_adr_o_i22 (.D(d_adr_o_31__N_2278[22]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[22] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i22.GSR = "ENABLED";
    FD1P3DX d_adr_o_i23 (.D(d_adr_o_31__N_2278[23]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[23] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i23.GSR = "ENABLED";
    FD1P3DX d_adr_o_i24 (.D(d_adr_o_31__N_2278[24]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[24] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i24.GSR = "ENABLED";
    FD1P3DX d_adr_o_i25 (.D(\d_adr_o_31__N_2278[25] ), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[25] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i25.GSR = "ENABLED";
    FD1P3DX d_adr_o_i26 (.D(d_adr_o_31__N_2278[26]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[26] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i26.GSR = "ENABLED";
    FD1P3DX d_adr_o_i27 (.D(\d_adr_o_31__N_2278[27] ), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[27] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i27.GSR = "ENABLED";
    FD1P3DX d_adr_o_i28 (.D(d_adr_o_31__N_2278[28]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[28] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i28.GSR = "ENABLED";
    FD1P3DX d_adr_o_i29 (.D(d_adr_o_31__N_2278[29]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[29] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i29.GSR = "ENABLED";
    FD1P3DX d_adr_o_i30 (.D(d_adr_o_31__N_2278[30]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[30] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i30.GSR = "ENABLED";
    FD1P3DX d_adr_o_i31 (.D(d_adr_o_31__N_2278[31]), .SP(REF_CLK_c_enable_1270), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32D_ADR_O[31] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i31.GSR = "ENABLED";
    FD1P3DX byte_enable_m_i0_i1 (.D(byte_enable_x[1]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(byte_enable_m[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam byte_enable_m_i0_i1.GSR = "ENABLED";
    FD1P3DX byte_enable_m_i0_i2 (.D(byte_enable_x[2]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(byte_enable_m[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam byte_enable_m_i0_i2.GSR = "ENABLED";
    FD1P3DX byte_enable_m_i0_i3 (.D(byte_enable_x[3]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(byte_enable_m[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam byte_enable_m_i0_i3.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i1 (.D(store_data_x[1]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i1.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i2 (.D(store_data_x[2]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i2.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i3 (.D(store_data_x[3]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i3.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i4 (.D(store_data_x[4]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i4.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i5 (.D(store_data_x[5]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i5.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i6 (.D(store_data_x[6]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i6.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i7 (.D(store_data_x[7]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i7.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i8 (.D(store_data_x[8]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i8.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i9 (.D(store_data_x[9]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i9.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i10 (.D(store_data_x[10]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i10.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i11 (.D(store_data_x[11]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i11.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i12 (.D(store_data_x[12]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i12.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i13 (.D(store_data_x[13]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i13.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i14 (.D(store_data_x[14]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i14.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i15 (.D(store_data_x[15]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i15.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i16 (.D(store_data_x[16]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i16.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i17 (.D(store_data_x[17]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i17.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i18 (.D(store_data_x[18]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i18.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i19 (.D(store_data_x[19]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i19.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i20 (.D(store_data_x[20]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i20.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i21 (.D(store_data_x[21]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i21.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i22 (.D(store_data_x[22]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i22.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i23 (.D(store_data_x[23]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i23.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i24 (.D(store_data_x[24]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i24.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i25 (.D(store_data_x[25]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i25.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i26 (.D(store_data_x[26]), .SP(REF_CLK_c_enable_1299), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i26.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i27 (.D(store_data_x[27]), .SP(REF_CLK_c_enable_1304), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i27.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i28 (.D(store_data_x[28]), .SP(REF_CLK_c_enable_1304), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i28.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i29 (.D(store_data_x[29]), .SP(REF_CLK_c_enable_1304), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i29.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i30 (.D(store_data_x[30]), .SP(REF_CLK_c_enable_1304), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i30.GSR = "ENABLED";
    FD1P3DX store_data_m_i0_i31 (.D(store_data_x[31]), .SP(REF_CLK_c_enable_1304), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(store_data_m[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i31.GSR = "ENABLED";
    FD1S3DX size_w_i1 (.D(size_m[1]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(size_w_c[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam size_w_i1.GSR = "ENABLED";
    FD1S3DX data_w_i1 (.D(data_m[1]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(data_w[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i1.GSR = "ENABLED";
    FD1S3DX data_w_i2 (.D(data_m[2]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(data_w[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i2.GSR = "ENABLED";
    FD1S3DX data_w_i3 (.D(data_m[3]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(data_w[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i3.GSR = "ENABLED";
    FD1S3DX data_w_i4 (.D(data_m[4]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(data_w[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i4.GSR = "ENABLED";
    FD1S3DX data_w_i5 (.D(data_m[5]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(data_w[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i5.GSR = "ENABLED";
    FD1S3DX data_w_i6 (.D(data_m[6]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(data_w[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i6.GSR = "ENABLED";
    FD1S3DX data_w_i7 (.D(data_m[7]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(data_w[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i7.GSR = "ENABLED";
    FD1S3DX data_w_i8 (.D(data_m[8]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\data_w[8] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i8.GSR = "ENABLED";
    FD1S3DX data_w_i9 (.D(data_m[9]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\data_w[9] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i9.GSR = "ENABLED";
    FD1S3DX data_w_i10 (.D(data_m[10]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\data_w[10] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i10.GSR = "ENABLED";
    FD1S3DX data_w_i11 (.D(data_m[11]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\data_w[11] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i11.GSR = "ENABLED";
    FD1S3DX data_w_i12 (.D(data_m[12]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\data_w[12] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i12.GSR = "ENABLED";
    FD1S3DX data_w_i13 (.D(data_m[13]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\data_w[13] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i13.GSR = "ENABLED";
    FD1S3DX data_w_i14 (.D(data_m[14]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\data_w[14] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i14.GSR = "ENABLED";
    FD1S3DX data_w_i15 (.D(data_m[15]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\data_w[15] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i15.GSR = "ENABLED";
    FD1S3DX data_w_i16 (.D(data_m[16]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(data_w[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i16.GSR = "ENABLED";
    FD1S3DX data_w_i17 (.D(data_m[17]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(data_w[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i17.GSR = "ENABLED";
    FD1S3DX data_w_i18 (.D(data_m[18]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(data_w[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i18.GSR = "ENABLED";
    FD1S3DX data_w_i19 (.D(data_m[19]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(data_w[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i19.GSR = "ENABLED";
    FD1S3DX data_w_i20 (.D(data_m[20]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(data_w[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i20.GSR = "ENABLED";
    FD1S3DX data_w_i21 (.D(data_m[21]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(data_w[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i21.GSR = "ENABLED";
    FD1S3DX data_w_i22 (.D(data_m[22]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(data_w[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i22.GSR = "ENABLED";
    FD1S3DX data_w_i23 (.D(data_m[23]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(data_w[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i23.GSR = "ENABLED";
    FD1S3DX data_w_i24 (.D(data_m[24]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\data_w[24] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i24.GSR = "ENABLED";
    FD1S3DX data_w_i25 (.D(data_m[25]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\data_w[25] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i25.GSR = "ENABLED";
    FD1S3DX data_w_i26 (.D(data_m[26]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\data_w[26] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i26.GSR = "ENABLED";
    FD1S3DX data_w_i27 (.D(data_m[27]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\data_w[27] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i27.GSR = "ENABLED";
    FD1S3DX data_w_i28 (.D(data_m[28]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\data_w[28] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i28.GSR = "ENABLED";
    FD1S3DX data_w_i29 (.D(data_m[29]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\data_w[29] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i29.GSR = "ENABLED";
    FD1S3DX data_w_i30 (.D(data_m[30]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\data_w[30] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i30.GSR = "ENABLED";
    FD1S3DX data_w_i31 (.D(data_m[31]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\data_w[31] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i31.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut_4_lut (.A(size_w_c[1]), .B(\operand_w[0] ), .C(data_w[23]), 
         .D(\data_w[31] ), .Z(n23_adj_6069)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_2_lut_4_lut_4_lut.init = 16'h5140;
    LUT4 i53_4_lut_4_lut (.A(size_w_c[1]), .B(\data_w[13] ), .C(\operand_w[0] ), 
         .D(data_w[5]), .Z(n28_adj_6076)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_4_lut.init = 16'hf404;
    LUT4 i53_4_lut_4_lut_adj_483 (.A(size_w_c[1]), .B(\data_w[11] ), .C(\operand_w[0] ), 
         .D(data_w[3]), .Z(n28_adj_6064)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_4_lut_adj_483.init = 16'hf404;
    LUT4 i1_4_lut_4_lut_adj_484 (.A(size_w_c[1]), .B(\operand_w[0] ), .C(data_w[21]), 
         .D(\data_w[29] ), .Z(n23_adj_6075)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_484.init = 16'h5140;
    LUT4 i1_4_lut_4_lut_adj_485 (.A(size_w_c[1]), .B(\operand_w[0] ), .C(data_w[19]), 
         .D(\data_w[27] ), .Z(n23_adj_6063)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_485.init = 16'h5140;
    LUT4 i53_4_lut_4_lut_adj_486 (.A(size_w_c[1]), .B(\data_w[12] ), .C(\operand_w[0] ), 
         .D(data_w[4]), .Z(n28_adj_6073)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_4_lut_adj_486.init = 16'hf404;
    LUT4 i53_4_lut_4_lut_adj_487 (.A(size_w_c[1]), .B(\data_w[10] ), .C(\operand_w[0] ), 
         .D(data_w[2]), .Z(n28_adj_6061)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_4_lut_adj_487.init = 16'hf404;
    LUT4 i1_4_lut_4_lut_adj_488 (.A(size_w_c[1]), .B(\operand_w[0] ), .C(data_w[20]), 
         .D(\data_w[28] ), .Z(n23_adj_6072)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_488.init = 16'h5140;
    LUT4 i1_4_lut_4_lut_adj_489 (.A(size_w_c[1]), .B(\operand_w[0] ), .C(data_w[18]), 
         .D(\data_w[26] ), .Z(n23_adj_6060)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_489.init = 16'h5140;
    LUT4 i53_4_lut_4_lut_adj_490 (.A(size_w_c[1]), .B(\data_w[15] ), .C(\operand_w[0] ), 
         .D(data_w[7]), .Z(n28_adj_6070)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_4_lut_adj_490.init = 16'hf404;
    LUT4 i53_4_lut_4_lut_adj_491 (.A(size_w_c[1]), .B(\data_w[9] ), .C(\operand_w[0] ), 
         .D(data_w[1]), .Z(n28_adj_6058)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_4_lut_adj_491.init = 16'hf404;
    LUT4 i1_4_lut_4_lut_adj_492 (.A(size_w_c[1]), .B(\operand_w[0] ), .C(data_w[17]), 
         .D(\data_w[25] ), .Z(n23_adj_6057)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_492.init = 16'h5140;
    LUT4 i53_4_lut_4_lut_adj_493 (.A(size_w_c[1]), .B(\data_w[14] ), .C(\operand_w[0] ), 
         .D(data_w[6]), .Z(n28_adj_6067)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_4_lut_adj_493.init = 16'hf404;
    LUT4 i53_4_lut_4_lut_adj_494 (.A(size_w_c[1]), .B(\data_w[8] ), .C(\operand_w[0] ), 
         .D(data_w[0]), .Z(n28)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_4_lut_adj_494.init = 16'hf404;
    LUT4 i1_4_lut_4_lut_adj_495 (.A(size_w_c[1]), .B(\operand_w[0] ), .C(data_w[22]), 
         .D(\data_w[30] ), .Z(n23_adj_6066)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_495.init = 16'h5140;
    LUT4 i1_4_lut_4_lut_adj_496 (.A(size_w_c[1]), .B(\operand_w[0] ), .C(data_w[16]), 
         .D(\data_w[24] ), .Z(n23)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_496.init = 16'h5140;
    LUT4 dcache_refilling_I_0_219_3_lut_rep_982 (.A(dcache_refilling), .B(\LM32D_ADR_O[2] ), 
         .C(\next_cycle_type[2] ), .Z(n41387)) /* synthesis lut_function=(!((B (C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(655[21:64])
    defparam dcache_refilling_I_0_219_3_lut_rep_982.init = 16'h2a2a;
    LUT4 i1_2_lut_3_lut (.A(dcache_refilling), .B(\LM32D_ADR_O[2] ), .C(\next_cycle_type[2] ), 
         .Z(n32298)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(655[21:64])
    defparam i1_2_lut_3_lut.init = 16'h0808;
    LUT4 i5092_4_lut_then_4_lut (.A(sign_extend_w), .B(data_w[7]), .C(\data_w[15] ), 
         .D(\operand_w[0] ), .Z(n41490)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i5092_4_lut_then_4_lut.init = 16'h88a0;
    LUT4 i5092_4_lut_else_4_lut (.A(sign_extend_w), .B(data_w[23]), .C(\data_w[31] ), 
         .D(\operand_w[0] ), .Z(n41489)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i5092_4_lut_else_4_lut.init = 16'h88a0;
    LUT4 i15373_2_lut (.A(dcache_refill_request), .B(LM32D_CYC_O), .Z(n20639)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i15373_2_lut.init = 16'heeee;
    LUT4 i3305_4_lut (.A(\LM32D_ADR_O[2] ), .B(n41380), .C(locked_N_493), 
         .D(n41387), .Z(n3722[0])) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(658[68:115])
    defparam i3305_4_lut.init = 16'h6aaa;
    LUT4 i3313_4_lut (.A(\next_cycle_type[2] ), .B(n32298), .C(locked_N_493), 
         .D(n41380), .Z(n3722[1])) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(658[68:115])
    defparam i3313_4_lut.init = 16'h6aaa;
    LUT4 i15107_2_lut (.A(operand_m[1]), .B(dcache_refill_request), .Z(d_adr_o_31__N_2278[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam i15107_2_lut.init = 16'h2222;
    LUT4 mux_99_i5_3_lut (.A(operand_m[4]), .B(dcache_refill_address[4]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i5_3_lut.init = 16'hcaca;
    LUT4 mux_99_i7_3_lut (.A(operand_m[6]), .B(dcache_refill_address[6]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i7_3_lut.init = 16'hcaca;
    LUT4 mux_99_i8_3_lut (.A(operand_m[7]), .B(dcache_refill_address[7]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i8_3_lut.init = 16'hcaca;
    LUT4 mux_99_i9_3_lut (.A(operand_m[8]), .B(dcache_refill_address[8]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i9_3_lut.init = 16'hcaca;
    LUT4 mux_99_i12_3_lut (.A(operand_m[11]), .B(dcache_refill_address[11]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i12_3_lut.init = 16'hcaca;
    LUT4 mux_99_i13_3_lut (.A(operand_m[12]), .B(dcache_refill_address[12]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i13_3_lut.init = 16'hcaca;
    LUT4 mux_99_i14_3_lut (.A(operand_m[13]), .B(dcache_refill_address[13]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i14_3_lut.init = 16'hcaca;
    LUT4 mux_99_i15_3_lut (.A(operand_m[14]), .B(dcache_refill_address[14]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i15_3_lut.init = 16'hcaca;
    LUT4 mux_99_i16_3_lut (.A(operand_m[15]), .B(dcache_refill_address[15]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i16_3_lut.init = 16'hcaca;
    LUT4 mux_99_i17_3_lut (.A(operand_m[16]), .B(dcache_refill_address[16]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i17_3_lut.init = 16'hcaca;
    LUT4 mux_99_i18_3_lut (.A(operand_m[17]), .B(dcache_refill_address[17]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i18_3_lut.init = 16'hcaca;
    LUT4 mux_99_i19_3_lut (.A(operand_m[18]), .B(dcache_refill_address[18]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i19_3_lut.init = 16'hcaca;
    LUT4 mux_99_i20_3_lut (.A(operand_m[19]), .B(dcache_refill_address[19]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i20_3_lut.init = 16'hcaca;
    LUT4 mux_99_i21_3_lut (.A(operand_m[20]), .B(dcache_refill_address[20]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i21_3_lut.init = 16'hcaca;
    LUT4 mux_99_i22_3_lut (.A(operand_m[21]), .B(dcache_refill_address[21]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i22_3_lut.init = 16'hcaca;
    LUT4 mux_99_i23_3_lut (.A(operand_m[22]), .B(dcache_refill_address[22]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i23_3_lut.init = 16'hcaca;
    LUT4 mux_99_i24_3_lut (.A(operand_m[23]), .B(dcache_refill_address[23]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i24_3_lut.init = 16'hcaca;
    LUT4 mux_99_i25_3_lut (.A(operand_m[24]), .B(dcache_refill_address[24]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i25_3_lut.init = 16'hcaca;
    LUT4 mux_99_i27_3_lut (.A(operand_m[26]), .B(dcache_refill_address[26]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i27_3_lut.init = 16'hcaca;
    LUT4 mux_99_i29_3_lut (.A(operand_m[28]), .B(dcache_refill_address[28]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i29_3_lut.init = 16'hcaca;
    LUT4 mux_99_i30_3_lut (.A(operand_m[29]), .B(dcache_refill_address[29]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i30_3_lut.init = 16'hcaca;
    LUT4 mux_99_i31_3_lut (.A(operand_m[30]), .B(dcache_refill_address[30]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i31_3_lut.init = 16'hcaca;
    LUT4 mux_99_i32_3_lut (.A(operand_m[31]), .B(dcache_refill_address[31]), 
         .C(dcache_refill_request), .Z(d_adr_o_31__N_2278[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam mux_99_i32_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut (.A(size_x[0]), .B(size_x[1]), .C(\adder_result_x[1] ), 
         .Z(n20800)) /* synthesis lut_function=(A ((C)+!B)+!A !(B)) */ ;
    defparam i1_3_lut.init = 16'hb3b3;
    LUT4 i14633_3_lut_4_lut (.A(n41215), .B(n41217), .C(dcache_refill_request), 
         .D(byte_enable_m[0]), .Z(d_sel_o_3__N_2358[0])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(718[18] 732[16])
    defparam i14633_3_lut_4_lut.init = 16'hfef0;
    LUT4 i15110_3_lut_4_lut (.A(n41215), .B(n41217), .C(dcache_refill_request), 
         .D(byte_enable_m[1]), .Z(d_sel_o_3__N_2358[1])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(718[18] 732[16])
    defparam i15110_3_lut_4_lut.init = 16'hfef0;
    LUT4 i15111_3_lut_4_lut (.A(n41215), .B(n41217), .C(dcache_refill_request), 
         .D(byte_enable_m[2]), .Z(d_sel_o_3__N_2358[2])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(718[18] 732[16])
    defparam i15111_3_lut_4_lut.init = 16'hfef0;
    LUT4 i15112_3_lut_4_lut (.A(n41215), .B(n41217), .C(dcache_refill_request), 
         .D(byte_enable_m[3]), .Z(d_sel_o_3__N_2358[3])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(718[18] 732[16])
    defparam i15112_3_lut_4_lut.init = 16'hfef0;
    LUT4 i2_2_lut_3_lut_4_lut (.A(n41215), .B(n41217), .C(LM32D_CYC_O), 
         .D(dcache_refill_request), .Z(REF_CLK_c_enable_1242)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(718[18] 732[16])
    defparam i2_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n41215), .B(n41217), .C(LM32D_CYC_O), 
         .D(dcache_refill_request), .Z(REF_CLK_c_enable_1270)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(718[18] 732[16])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0f0e;
    LUT4 size_x_1__I_0_192_Mux_24_i2_3_lut (.A(store_operand_x[24]), .B(store_operand_x[8]), 
         .C(size_x[0]), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_24_i2_3_lut.init = 16'hcaca;
    LUT4 size_x_1__I_0_192_Mux_25_i2_3_lut (.A(store_operand_x[25]), .B(store_operand_x[9]), 
         .C(size_x[0]), .Z(n2_adj_6084)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_25_i2_3_lut.init = 16'hcaca;
    LUT4 size_x_1__I_0_192_Mux_26_i2_3_lut (.A(store_operand_x[26]), .B(store_operand_x[10]), 
         .C(size_x[0]), .Z(n2_adj_6085)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_26_i2_3_lut.init = 16'hcaca;
    LUT4 size_x_1__I_0_192_Mux_27_i2_3_lut (.A(store_operand_x[27]), .B(store_operand_x[11]), 
         .C(size_x[0]), .Z(n2_adj_6086)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_27_i2_3_lut.init = 16'hcaca;
    LUT4 size_x_1__I_0_192_Mux_28_i2_3_lut (.A(store_operand_x[28]), .B(store_operand_x[12]), 
         .C(size_x[0]), .Z(n2_adj_6087)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_28_i2_3_lut.init = 16'hcaca;
    LUT4 size_x_1__I_0_192_Mux_29_i2_3_lut (.A(store_operand_x[29]), .B(store_operand_x[13]), 
         .C(size_x[0]), .Z(n2_adj_6088)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_29_i2_3_lut.init = 16'hcaca;
    LUT4 size_x_1__I_0_192_Mux_30_i2_3_lut (.A(store_operand_x[30]), .B(store_operand_x[14]), 
         .C(size_x[0]), .Z(n2_adj_6089)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_30_i2_3_lut.init = 16'hcaca;
    LUT4 size_x_1__I_0_192_Mux_31_i2_3_lut (.A(store_operand_x[31]), .B(store_operand_x[15]), 
         .C(size_x[0]), .Z(n2_adj_6090)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_31_i2_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i2_3_lut (.A(dcache_data_m[1]), .B(wb_data_m[1]), 
         .C(wb_select_m), .Z(data_m[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i3_3_lut (.A(dcache_data_m[2]), .B(wb_data_m[2]), 
         .C(wb_select_m), .Z(data_m[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i4_3_lut (.A(dcache_data_m[3]), .B(wb_data_m[3]), 
         .C(wb_select_m), .Z(data_m[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i5_3_lut (.A(dcache_data_m[4]), .B(wb_data_m[4]), 
         .C(wb_select_m), .Z(data_m[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i6_3_lut (.A(dcache_data_m[5]), .B(wb_data_m[5]), 
         .C(wb_select_m), .Z(data_m[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i7_3_lut (.A(dcache_data_m[6]), .B(wb_data_m[6]), 
         .C(wb_select_m), .Z(data_m[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i8_3_lut (.A(dcache_data_m[7]), .B(wb_data_m[7]), 
         .C(wb_select_m), .Z(data_m[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i9_3_lut (.A(n6416[0]), .B(wb_data_m[8]), 
         .C(wb_select_m), .Z(data_m[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i10_3_lut (.A(n6416[1]), .B(wb_data_m[9]), 
         .C(wb_select_m), .Z(data_m[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i11_3_lut (.A(n6416[2]), .B(wb_data_m[10]), 
         .C(wb_select_m), .Z(data_m[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i12_3_lut (.A(n6416[3]), .B(wb_data_m[11]), 
         .C(wb_select_m), .Z(data_m[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i13_3_lut (.A(n6416[4]), .B(wb_data_m[12]), 
         .C(wb_select_m), .Z(data_m[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i13_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i14_3_lut (.A(n6416[5]), .B(wb_data_m[13]), 
         .C(wb_select_m), .Z(data_m[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i14_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i15_3_lut (.A(n6416[6]), .B(wb_data_m[14]), 
         .C(wb_select_m), .Z(data_m[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i15_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i16_3_lut (.A(n6416[7]), .B(wb_data_m[15]), 
         .C(wb_select_m), .Z(data_m[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i16_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i17_3_lut (.A(n6417[0]), .B(wb_data_m[16]), 
         .C(wb_select_m), .Z(data_m[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i17_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i18_3_lut (.A(n6417[1]), .B(wb_data_m[17]), 
         .C(wb_select_m), .Z(data_m[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i18_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i19_3_lut (.A(n6417[2]), .B(wb_data_m[18]), 
         .C(wb_select_m), .Z(data_m[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i19_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i20_3_lut (.A(n6417[3]), .B(wb_data_m[19]), 
         .C(wb_select_m), .Z(data_m[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i20_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_adj_497 (.A(size_x[1]), .B(size_x[0]), .C(\adder_result_x[1] ), 
         .Z(n9_c)) /* synthesis lut_function=(A ((C)+!B)) */ ;
    defparam i1_3_lut_adj_497.init = 16'ha2a2;
    LUT4 kill_m_I_0_2_lut_rep_987 (.A(dcache_refill_request), .B(exception_m), 
         .Z(n41392)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(741[13:56])
    defparam kill_m_I_0_2_lut_rep_987.init = 16'heeee;
    LUT4 i30535_2_lut_3_lut (.A(dcache_refill_request), .B(exception_m), 
         .C(dcache_select_x), .Z(n35694)) /* synthesis lut_function=(A+(B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(741[13:56])
    defparam i30535_2_lut_3_lut.init = 16'hfefe;
    LUT4 dcache_data_m_31__I_0_i21_3_lut (.A(n6417[4]), .B(wb_data_m[20]), 
         .C(wb_select_m), .Z(data_m[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i21_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i22_3_lut (.A(n6417[5]), .B(wb_data_m[21]), 
         .C(wb_select_m), .Z(data_m[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i22_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i23_3_lut (.A(n6417[6]), .B(wb_data_m[22]), 
         .C(wb_select_m), .Z(data_m[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i23_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i24_3_lut (.A(n6417[7]), .B(wb_data_m[23]), 
         .C(wb_select_m), .Z(data_m[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i24_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i25_3_lut (.A(n6418[0]), .B(wb_data_m[24]), 
         .C(wb_select_m), .Z(data_m[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i25_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i26_3_lut (.A(n6418[1]), .B(wb_data_m[25]), 
         .C(wb_select_m), .Z(data_m[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i26_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i27_3_lut (.A(n6418[2]), .B(wb_data_m[26]), 
         .C(wb_select_m), .Z(data_m[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i27_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i28_3_lut (.A(n6418[3]), .B(wb_data_m[27]), 
         .C(wb_select_m), .Z(data_m[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i28_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i1_3_lut (.A(dcache_data_m[0]), .B(wb_data_m[0]), 
         .C(wb_select_m), .Z(data_m[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i29_3_lut (.A(n6418[4]), .B(wb_data_m[28]), 
         .C(wb_select_m), .Z(data_m[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i29_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i30_3_lut (.A(n6418[5]), .B(wb_data_m[29]), 
         .C(wb_select_m), .Z(data_m[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i30_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i31_3_lut (.A(n6418[6]), .B(wb_data_m[30]), 
         .C(wb_select_m), .Z(data_m[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i31_3_lut.init = 16'hcaca;
    LUT4 dcache_data_m_31__I_0_i32_3_lut (.A(n6418[7]), .B(wb_data_m[31]), 
         .C(wb_select_m), .Z(data_m[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(538[20] 540[35])
    defparam dcache_data_m_31__I_0_i32_3_lut.init = 16'hcaca;
    LUT4 i15381_2_lut_3_lut (.A(size_x[0]), .B(size_x[1]), .C(store_operand_x[3]), 
         .Z(store_data_x[3])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam i15381_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i15383_2_lut_3_lut (.A(size_x[0]), .B(size_x[1]), .C(store_operand_x[1]), 
         .Z(store_data_x[1])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam i15383_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i1_4_lut_adj_498 (.A(n34978), .B(n41215), .C(n41217), .D(n20639), 
         .Z(REF_CLK_c_enable_193)) /* synthesis lut_function=(A+!((C+(D))+!B)) */ ;
    defparam i1_4_lut_adj_498.init = 16'haaae;
    LUT4 i1_4_lut_adj_499 (.A(n41232), .B(n41392), .C(n30070), .D(n35745), 
         .Z(n34978)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut_adj_499.init = 16'hccec;
    LUT4 i1_4_lut_adj_500 (.A(n41232), .B(n30070), .C(n41233), .D(n35694), 
         .Z(n31463)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_500.init = 16'h0008;
    LUT4 i15368_2_lut_3_lut (.A(size_x[0]), .B(size_x[1]), .C(store_operand_x[0]), 
         .Z(store_data_x[0])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam i15368_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i15382_2_lut_3_lut (.A(size_x[0]), .B(size_x[1]), .C(store_operand_x[2]), 
         .Z(store_data_x[2])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam i15382_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i15380_2_lut_3_lut (.A(size_x[0]), .B(size_x[1]), .C(store_operand_x[4]), 
         .Z(store_data_x[4])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam i15380_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i15379_2_lut_3_lut (.A(size_x[0]), .B(size_x[1]), .C(store_operand_x[5]), 
         .Z(store_data_x[5])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam i15379_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i15378_2_lut_3_lut (.A(size_x[0]), .B(size_x[1]), .C(store_operand_x[6]), 
         .Z(store_data_x[6])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam i15378_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i15377_2_lut_3_lut (.A(size_x[0]), .B(size_x[1]), .C(store_operand_x[7]), 
         .Z(store_data_x[7])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam i15377_2_lut_3_lut.init = 16'hd0d0;
    LUT4 dcache_select_x_I_0_1_lut (.A(dcache_select_x), .Z(dcache_select_x_N_2440)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(436[28:44])
    defparam dcache_select_x_I_0_1_lut.init = 16'h5555;
    LUT4 i23_3_lut (.A(n11), .B(n9), .C(LM32D_CYC_O), .Z(REF_CLK_c_enable_398)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23_3_lut.init = 16'hcaca;
    LUT4 i7014_3_lut (.A(n11), .B(n9), .C(LM32D_CYC_O), .Z(n12384)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam i7014_3_lut.init = 16'h3a3a;
    LUT4 i1_4_lut_4_lut_adj_501 (.A(data_w[16]), .B(data_w[0]), .C(\operand_w[1] ), 
         .D(size_w[0]), .Z(n25_adj_6092)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_501.init = 16'hcacc;
    LUT4 i1_4_lut_4_lut_adj_502 (.A(size_w[0]), .B(n31_adj_6068), .C(n25_adj_6082), 
         .D(size_w_c[1]), .Z(\load_data_w[6] )) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_502.init = 16'hf444;
    LUT4 n33_bdd_3_lut_34331_4_lut_4_lut (.A(size_w[0]), .B(n41144), .C(size_w_c[1]), 
         .D(n35), .Z(n41145)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam n33_bdd_3_lut_34331_4_lut_4_lut.init = 16'hc5c0;
    LUT4 n33_bdd_3_lut_34346_4_lut_4_lut (.A(size_w[0]), .B(n41156), .C(size_w_c[1]), 
         .D(n35), .Z(n41157)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam n33_bdd_3_lut_34346_4_lut_4_lut.init = 16'hc5c0;
    LUT4 n33_bdd_3_lut_34326_4_lut_4_lut (.A(size_w[0]), .B(n41140), .C(size_w_c[1]), 
         .D(n35), .Z(n41141)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam n33_bdd_3_lut_34326_4_lut_4_lut.init = 16'hc5c0;
    LUT4 n33_bdd_3_lut_4_lut_4_lut (.A(size_w[0]), .B(n41164), .C(size_w_c[1]), 
         .D(n35), .Z(n41165)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam n33_bdd_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 n33_bdd_3_lut_34351_4_lut_4_lut (.A(size_w[0]), .B(n41160), .C(size_w_c[1]), 
         .D(n35), .Z(n41161)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam n33_bdd_3_lut_34351_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i1_4_lut_4_lut_adj_503 (.A(size_w[0]), .B(n31_adj_6071), .C(n25_adj_6083), 
         .D(size_w_c[1]), .Z(\load_data_w[7] )) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_503.init = 16'hf444;
    LUT4 i1_4_lut_4_lut_adj_504 (.A(size_w[0]), .B(n31_adj_6077), .C(n25_adj_6081), 
         .D(size_w_c[1]), .Z(\load_data_w[5] )) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_504.init = 16'hf444;
    LUT4 i1_4_lut_4_lut_adj_505 (.A(size_w[0]), .B(n31_adj_6074), .C(n25_adj_6080), 
         .D(size_w_c[1]), .Z(\load_data_w[4] )) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_505.init = 16'hf444;
    LUT4 n33_bdd_3_lut_34336_4_lut_4_lut (.A(size_w[0]), .B(n41148), .C(size_w_c[1]), 
         .D(n35), .Z(n41149)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam n33_bdd_3_lut_34336_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i1_4_lut_4_lut_adj_506 (.A(size_w[0]), .B(n31_adj_6065), .C(n25_adj_6079), 
         .D(size_w_c[1]), .Z(\load_data_w[3] )) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_506.init = 16'hf444;
    LUT4 n33_bdd_3_lut_34341_4_lut_4_lut (.A(size_w[0]), .B(n41152), .C(size_w_c[1]), 
         .D(n35), .Z(n41153)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam n33_bdd_3_lut_34341_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i1_4_lut_4_lut_adj_507 (.A(size_w[0]), .B(n31_adj_6062), .C(n25_adj_6078), 
         .D(size_w_c[1]), .Z(\load_data_w[2] )) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_507.init = 16'hf444;
    LUT4 n33_bdd_3_lut_34321_4_lut_4_lut (.A(size_w[0]), .B(n41136), .C(size_w_c[1]), 
         .D(n35), .Z(n41137)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam n33_bdd_3_lut_34321_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i1_4_lut_4_lut_adj_508 (.A(size_w[0]), .B(n31_adj_6059), .C(n25), 
         .D(size_w_c[1]), .Z(\load_data_w[1] )) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_508.init = 16'hf444;
    LUT4 i1_4_lut_4_lut_adj_509 (.A(size_w[0]), .B(n31), .C(n25_adj_6092), 
         .D(size_w_c[1]), .Z(\load_data_w[0] )) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_509.init = 16'hf444;
    LUT4 i1_2_lut_rep_1030 (.A(dcache_refill_request), .B(icache_refill_request), 
         .Z(n41435)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam i1_2_lut_rep_1030.init = 16'heeee;
    LUT4 i1_2_lut_rep_798_3_lut (.A(dcache_refill_request), .B(icache_refill_request), 
         .C(branch_taken_m), .Z(n41203)) /* synthesis lut_function=(A+(B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam i1_2_lut_rep_798_3_lut.init = 16'hfefe;
    LUT4 valid_d_I_0_2_lut_3_lut_4_lut (.A(dcache_refill_request), .B(icache_refill_request), 
         .C(valid_d), .D(branch_taken_m), .Z(q_d)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam valid_d_I_0_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_3_lut_4_lut_adj_510 (.A(dcache_refill_request), .B(icache_refill_request), 
         .C(valid_d), .D(branch_taken_m), .Z(n32652)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(699[18] 732[16])
    defparam i1_3_lut_4_lut_adj_510.init = 16'hffef;
    LUT4 size_x_1__I_0_192_Mux_15_i3_3_lut_4_lut (.A(store_operand_x[7]), 
         .B(size_x[0]), .C(size_x[1]), .D(store_operand_x[15]), .Z(store_data_x[15])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_15_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_192_Mux_31_i3_3_lut_4_lut (.A(store_operand_x[7]), 
         .B(size_x[0]), .C(size_x[1]), .D(n2_adj_6090), .Z(store_data_x[31])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_31_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_192_Mux_14_i3_3_lut_4_lut (.A(store_operand_x[6]), 
         .B(size_x[0]), .C(size_x[1]), .D(store_operand_x[14]), .Z(store_data_x[14])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_14_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_192_Mux_30_i3_3_lut_4_lut (.A(store_operand_x[6]), 
         .B(size_x[0]), .C(size_x[1]), .D(n2_adj_6089), .Z(store_data_x[30])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_30_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_192_Mux_13_i3_3_lut_4_lut (.A(store_operand_x[5]), 
         .B(size_x[0]), .C(size_x[1]), .D(store_operand_x[13]), .Z(store_data_x[13])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_13_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_192_Mux_29_i3_3_lut_4_lut (.A(store_operand_x[5]), 
         .B(size_x[0]), .C(size_x[1]), .D(n2_adj_6088), .Z(store_data_x[29])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_29_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_192_Mux_12_i3_3_lut_4_lut (.A(store_operand_x[4]), 
         .B(size_x[0]), .C(size_x[1]), .D(store_operand_x[12]), .Z(store_data_x[12])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_12_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_192_Mux_28_i3_3_lut_4_lut (.A(store_operand_x[4]), 
         .B(size_x[0]), .C(size_x[1]), .D(n2_adj_6087), .Z(store_data_x[28])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_28_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_192_Mux_11_i3_3_lut_4_lut (.A(store_operand_x[3]), 
         .B(size_x[0]), .C(size_x[1]), .D(store_operand_x[11]), .Z(store_data_x[11])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_11_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_192_Mux_27_i3_3_lut_4_lut (.A(store_operand_x[3]), 
         .B(size_x[0]), .C(size_x[1]), .D(n2_adj_6086), .Z(store_data_x[27])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_27_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_192_Mux_10_i3_3_lut_4_lut (.A(store_operand_x[2]), 
         .B(size_x[0]), .C(size_x[1]), .D(store_operand_x[10]), .Z(store_data_x[10])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_10_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_192_Mux_26_i3_3_lut_4_lut (.A(store_operand_x[2]), 
         .B(size_x[0]), .C(size_x[1]), .D(n2_adj_6085), .Z(store_data_x[26])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_26_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_192_Mux_9_i3_3_lut_4_lut (.A(store_operand_x[1]), .B(size_x[0]), 
         .C(size_x[1]), .D(store_operand_x[9]), .Z(store_data_x[9])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_9_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_192_Mux_25_i3_3_lut_4_lut (.A(store_operand_x[1]), 
         .B(size_x[0]), .C(size_x[1]), .D(n2_adj_6084), .Z(store_data_x[25])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_25_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_192_Mux_8_i3_3_lut_4_lut (.A(store_operand_x[0]), .B(size_x[0]), 
         .C(size_x[1]), .D(store_operand_x[8]), .Z(store_data_x[8])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_8_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_192_Mux_24_i3_3_lut_4_lut (.A(store_operand_x[0]), 
         .B(size_x[0]), .C(size_x[1]), .D(n2), .Z(store_data_x[24])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_192_Mux_24_i3_3_lut_4_lut.init = 16'hf202;
    PFUMX d_adr_o_31__I_0_i4 (.BLUT(\d_adr_o_31__N_2278[3] ), .ALUT(n3722[1]), 
          .C0(LM32D_CYC_O), .Z(d_adr_o_31__N_2149[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;
    PFUMX d_adr_o_31__I_0_i3 (.BLUT(\d_adr_o_31__N_2278[2] ), .ALUT(n3722[0]), 
          .C0(LM32D_CYC_O), .Z(d_adr_o_31__N_2149[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;
    \lm32_dcache(base_address=32'b0,limit=32'b01111111111111111)  dcache (.dcache_restart_request(dcache_restart_request), 
            .n45183(n45183), .state({state}), .REF_CLK_c(REF_CLK_c), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .flush_set({flush_set}), .flush_set_8__N_2513({flush_set_8__N_2513}), 
            .\dcache_refill_address[4] (dcache_refill_address[4]), .\operand_m[4] (operand_m[4]), 
            .dcache_refill_request(dcache_refill_request), .dcache_refilling(dcache_refilling), 
            .\dcache_refill_address[5] (\dcache_refill_address[5] ), .\operand_m[5] (operand_m[5]), 
            .\dcache_refill_address[6] (dcache_refill_address[6]), .\operand_m[6] (operand_m[6]), 
            .\dcache_refill_address[7] (dcache_refill_address[7]), .\operand_m[7] (operand_m[7]), 
            .\dcache_refill_address[8] (dcache_refill_address[8]), .\operand_m[8] (operand_m[8]), 
            .\dcache_refill_address[9] (\dcache_refill_address[9] ), .\operand_m[9] (operand_m[9]), 
            .\dcache_refill_address[10] (\dcache_refill_address[10] ), .\operand_m[10] (operand_m[10]), 
            .\dcache_refill_address[11] (dcache_refill_address[11]), .\operand_m[11] (operand_m[11]), 
            .\dcache_refill_address[12] (dcache_refill_address[12]), .\operand_m[12] (operand_m[12]), 
            .\dcache_refill_address[13] (dcache_refill_address[13]), .\operand_m[13] (operand_m[13]), 
            .\dcache_refill_address[14] (dcache_refill_address[14]), .\operand_m[14] (operand_m[14]), 
            .\dcache_refill_address[15] (dcache_refill_address[15]), .\operand_m[15] (operand_m[15]), 
            .\dcache_refill_address[16] (dcache_refill_address[16]), .\operand_m[16] (operand_m[16]), 
            .\dcache_refill_address[17] (dcache_refill_address[17]), .\operand_m[17] (operand_m[17]), 
            .\dcache_refill_address[18] (dcache_refill_address[18]), .\operand_m[18] (operand_m[18]), 
            .\dcache_refill_address[19] (dcache_refill_address[19]), .\operand_m[19] (operand_m[19]), 
            .\dcache_refill_address[20] (dcache_refill_address[20]), .\operand_m[20] (operand_m[20]), 
            .\dcache_refill_address[21] (dcache_refill_address[21]), .\operand_m[21] (operand_m[21]), 
            .\dcache_refill_address[22] (dcache_refill_address[22]), .\operand_m[22] (operand_m[22]), 
            .\dcache_refill_address[23] (dcache_refill_address[23]), .\operand_m[23] (operand_m[23]), 
            .\dcache_refill_address[24] (dcache_refill_address[24]), .\operand_m[24] (operand_m[24]), 
            .\dcache_refill_address[25] (\dcache_refill_address[25] ), .\operand_m[25] (operand_m[25]), 
            .\dcache_refill_address[26] (dcache_refill_address[26]), .\operand_m[26] (operand_m[26]), 
            .\dcache_refill_address[27] (\dcache_refill_address[27] ), .\operand_m[27] (operand_m[27]), 
            .\dcache_refill_address[28] (dcache_refill_address[28]), .\operand_m[28] (operand_m[28]), 
            .\dcache_refill_address[29] (dcache_refill_address[29]), .\operand_m[29] (operand_m[29]), 
            .\dcache_refill_address[30] (dcache_refill_address[30]), .\operand_m[30] (operand_m[30]), 
            .\dcache_refill_address[31] (dcache_refill_address[31]), .\operand_m[31] (operand_m[31]), 
            .store_data_m({store_data_m}), .wb_data_m({wb_data_m}), .n45171(n45171), 
            .n41284(n41284), .dcache_select_m(dcache_select_m), .n41435(n41435), 
            .icache_restart_request(icache_restart_request), .n19852(n19852), 
            .valid_a(valid_a), .n30107(n30107), .dcache_refill_ready(dcache_refill_ready), 
            .n41233(n41233), .\operand_m[2] (operand_m[2]), .\operand_m[3] (operand_m[3]), 
            .n9304(n9304), .\state[2]_adj_181 (\state[2]_adj_192 ), .n41187(n41187), 
            .n41196(n41196), .n41203(n41203), .n31996(n31996), .n45175(n45175), 
            .way_match_0__N_2007(way_match_0__N_2007), .valid_f(valid_f), 
            .\operand_m[0] (operand_m[0]), .\d_adr_o_31__N_2278[0] (d_adr_o_31__N_2278[0]), 
            .dflush_m(dflush_m), .branch_taken_m(branch_taken_m), .n41178(n41178), 
            .n36389(n36389), .n37914(n37914), .n37915(n37915), .n37919(n37919), 
            .n37917(n37917), .n37916(n37916), .n37918(n37918), .n41(n41), 
            .icache_refill_request(icache_refill_request), .restart_request_N_1998(restart_request_N_1998), 
            .n15(n15), .n41172(n41172), .n32278(n32278), .\tmem_write_address[1] (\tmem_write_address[1] ), 
            .\tmem_write_address[5] (\tmem_write_address[5] ), .\tmem_write_address[6] (\tmem_write_address[6] ), 
            .n7502({n7502}), .VCC_net(VCC_net), .GND_net(GND_net), .\genblk1.ra ({\genblk1.ra }), 
            .\dmem_write_address[3] (\dmem_write_address[3] ), .\dmem_write_address[7] (\dmem_write_address[7] ), 
            .\dmem_write_address[8] (\dmem_write_address[8] ), .n7388({n7388}), 
            .byte_enable_m({byte_enable_m}), .n7322({n7322}), .n7256({n7256}), 
            .n7204(n7204), .n7190({n7190}), .n7206(n7206), .n7208(n7208), 
            .\genblk1.ra_adj_191 ({\genblk1.ra_adj_202 }), .n6418({n6418}), 
            .n7224(n7224), .n7222(n7222), .n7220(n7220), .n6417({n6417}), 
            .n7356(n7356), .n7354(n7354), .n7352(n7352), .n7350(n7350), 
            .n7348(n7348), .n7346(n7346), .n7344(n7344), .n7342(n7342), 
            .n7340(n7340), .n7338(n7338), .n7336(n7336), .n7218(n7218), 
            .n7290(n7290), .n7288(n7288), .n7286(n7286), .n7284(n7284), 
            .n7216(n7216), .n7282(n7282), .n6416({n6416}), .n7280(n7280), 
            .n7278(n7278), .n7214(n7214), .n7276(n7276), .n7274(n7274), 
            .n7272(n7272), .n7212(n7212), .n7270(n7270), .n7210(n7210), 
            .dcache_data_m({dcache_data_m})) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(381[7] 404[6])
    
endmodule
//
// Verilog Description of module \lm32_dcache(base_address=32'b0,limit=32'b01111111111111111) 
//

module \lm32_dcache(base_address=32'b0,limit=32'b01111111111111111)  (dcache_restart_request, 
            n45183, state, REF_CLK_c, REF_CLK_c_enable_1606, flush_set, 
            flush_set_8__N_2513, \dcache_refill_address[4] , \operand_m[4] , 
            dcache_refill_request, dcache_refilling, \dcache_refill_address[5] , 
            \operand_m[5] , \dcache_refill_address[6] , \operand_m[6] , 
            \dcache_refill_address[7] , \operand_m[7] , \dcache_refill_address[8] , 
            \operand_m[8] , \dcache_refill_address[9] , \operand_m[9] , 
            \dcache_refill_address[10] , \operand_m[10] , \dcache_refill_address[11] , 
            \operand_m[11] , \dcache_refill_address[12] , \operand_m[12] , 
            \dcache_refill_address[13] , \operand_m[13] , \dcache_refill_address[14] , 
            \operand_m[14] , \dcache_refill_address[15] , \operand_m[15] , 
            \dcache_refill_address[16] , \operand_m[16] , \dcache_refill_address[17] , 
            \operand_m[17] , \dcache_refill_address[18] , \operand_m[18] , 
            \dcache_refill_address[19] , \operand_m[19] , \dcache_refill_address[20] , 
            \operand_m[20] , \dcache_refill_address[21] , \operand_m[21] , 
            \dcache_refill_address[22] , \operand_m[22] , \dcache_refill_address[23] , 
            \operand_m[23] , \dcache_refill_address[24] , \operand_m[24] , 
            \dcache_refill_address[25] , \operand_m[25] , \dcache_refill_address[26] , 
            \operand_m[26] , \dcache_refill_address[27] , \operand_m[27] , 
            \dcache_refill_address[28] , \operand_m[28] , \dcache_refill_address[29] , 
            \operand_m[29] , \dcache_refill_address[30] , \operand_m[30] , 
            \dcache_refill_address[31] , \operand_m[31] , store_data_m, 
            wb_data_m, n45171, n41284, dcache_select_m, n41435, icache_restart_request, 
            n19852, valid_a, n30107, dcache_refill_ready, n41233, 
            \operand_m[2] , \operand_m[3] , n9304, \state[2]_adj_181 , 
            n41187, n41196, n41203, n31996, n45175, way_match_0__N_2007, 
            valid_f, \operand_m[0] , \d_adr_o_31__N_2278[0] , dflush_m, 
            branch_taken_m, n41178, n36389, n37914, n37915, n37919, 
            n37917, n37916, n37918, n41, icache_refill_request, restart_request_N_1998, 
            n15, n41172, n32278, \tmem_write_address[1] , \tmem_write_address[5] , 
            \tmem_write_address[6] , n7502, VCC_net, GND_net, \genblk1.ra , 
            \dmem_write_address[3] , \dmem_write_address[7] , \dmem_write_address[8] , 
            n7388, byte_enable_m, n7322, n7256, n7204, n7190, n7206, 
            n7208, \genblk1.ra_adj_191 , n6418, n7224, n7222, n7220, 
            n6417, n7356, n7354, n7352, n7350, n7348, n7346, n7344, 
            n7342, n7340, n7338, n7336, n7218, n7290, n7288, n7286, 
            n7284, n7216, n7282, n6416, n7280, n7278, n7214, n7276, 
            n7274, n7272, n7212, n7270, n7210, dcache_data_m) /* synthesis syn_module_defined=1 */ ;
    output dcache_restart_request;
    input n45183;
    output [2:0]state;
    input REF_CLK_c;
    input REF_CLK_c_enable_1606;
    output [8:0]flush_set;
    input [8:0]flush_set_8__N_2513;
    output \dcache_refill_address[4] ;
    input \operand_m[4] ;
    output dcache_refill_request;
    output dcache_refilling;
    output \dcache_refill_address[5] ;
    input \operand_m[5] ;
    output \dcache_refill_address[6] ;
    input \operand_m[6] ;
    output \dcache_refill_address[7] ;
    input \operand_m[7] ;
    output \dcache_refill_address[8] ;
    input \operand_m[8] ;
    output \dcache_refill_address[9] ;
    input \operand_m[9] ;
    output \dcache_refill_address[10] ;
    input \operand_m[10] ;
    output \dcache_refill_address[11] ;
    input \operand_m[11] ;
    output \dcache_refill_address[12] ;
    input \operand_m[12] ;
    output \dcache_refill_address[13] ;
    input \operand_m[13] ;
    output \dcache_refill_address[14] ;
    input \operand_m[14] ;
    output \dcache_refill_address[15] ;
    input \operand_m[15] ;
    output \dcache_refill_address[16] ;
    input \operand_m[16] ;
    output \dcache_refill_address[17] ;
    input \operand_m[17] ;
    output \dcache_refill_address[18] ;
    input \operand_m[18] ;
    output \dcache_refill_address[19] ;
    input \operand_m[19] ;
    output \dcache_refill_address[20] ;
    input \operand_m[20] ;
    output \dcache_refill_address[21] ;
    input \operand_m[21] ;
    output \dcache_refill_address[22] ;
    input \operand_m[22] ;
    output \dcache_refill_address[23] ;
    input \operand_m[23] ;
    output \dcache_refill_address[24] ;
    input \operand_m[24] ;
    output \dcache_refill_address[25] ;
    input \operand_m[25] ;
    output \dcache_refill_address[26] ;
    input \operand_m[26] ;
    output \dcache_refill_address[27] ;
    input \operand_m[27] ;
    output \dcache_refill_address[28] ;
    input \operand_m[28] ;
    output \dcache_refill_address[29] ;
    input \operand_m[29] ;
    output \dcache_refill_address[30] ;
    input \operand_m[30] ;
    output \dcache_refill_address[31] ;
    input \operand_m[31] ;
    input [31:0]store_data_m;
    input [31:0]wb_data_m;
    input n45171;
    input n41284;
    input dcache_select_m;
    input n41435;
    input icache_restart_request;
    input n19852;
    output valid_a;
    input n30107;
    input dcache_refill_ready;
    input n41233;
    input \operand_m[2] ;
    input \operand_m[3] ;
    input n9304;
    input \state[2]_adj_181 ;
    input n41187;
    input n41196;
    input n41203;
    output n31996;
    input n45175;
    input way_match_0__N_2007;
    input valid_f;
    input \operand_m[0] ;
    output \d_adr_o_31__N_2278[0] ;
    input dflush_m;
    input branch_taken_m;
    output n41178;
    output n36389;
    output n37914;
    output n37915;
    output n37919;
    output n37917;
    output n37916;
    output n37918;
    input n41;
    input icache_refill_request;
    output restart_request_N_1998;
    input n15;
    output n41172;
    output n32278;
    input \tmem_write_address[1] ;
    input \tmem_write_address[5] ;
    input \tmem_write_address[6] ;
    input [8:0]n7502;
    input VCC_net;
    input GND_net;
    output [8:0]\genblk1.ra ;
    input \dmem_write_address[3] ;
    input \dmem_write_address[7] ;
    input \dmem_write_address[8] ;
    input [10:0]n7388;
    input [3:0]byte_enable_m;
    input [10:0]n7322;
    input [10:0]n7256;
    output n7204;
    input [10:0]n7190;
    output n7206;
    output n7208;
    output [10:0]\genblk1.ra_adj_191 ;
    output [7:0]n6418;
    output n7224;
    output n7222;
    output n7220;
    output [7:0]n6417;
    output n7356;
    output n7354;
    output n7352;
    output n7350;
    output n7348;
    output n7346;
    output n7344;
    output n7342;
    output n7340;
    output n7338;
    output n7336;
    output n7218;
    output n7290;
    output n7288;
    output n7286;
    output n7284;
    output n7216;
    output n7282;
    output [7:0]n6416;
    output n7280;
    output n7278;
    output n7214;
    output n7276;
    output n7274;
    output n7272;
    output n7212;
    output n7270;
    output n7210;
    output [7:0]dcache_data_m;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    
    wire n38909, n9244, REF_CLK_c_enable_1480;
    wire [3:2]refill_offset;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(193[32:45])
    wire [1:0]refill_offset_3__N_2489;
    
    wire refill_request_N_2565, restart_request_N_2560, n31551, n9248;
    wire [31:0]dmem_write_data;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(184[22:37])
    
    wire way_match_0__N_2572, miss;
    wire [3:0]way_valid;
    
    wire n4, n2, n3, n7540, n7541, n41218, n7536, n7537, n7538, 
        n7539, n9291;
    wire [10:0]dmem_write_address;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(182[31:49])
    wire [8:0]tmem_write_address;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(180[31:49])
    wire [0:0]way_tmem_we;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(171[26:37])
    
    wire n36, n31990, n4_adj_6029;
    wire [1:0]refill_offset_3__N_2557;
    
    wire n41176, n34780, n41320, n23436, n35822, n35824, n35512, 
        n31665, n35540, n35538, n38908;
    wire [3:0]tmem_write_data;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(183[26:41])
    
    wire n7426, n7428, n7430, n7432, n7434, n7436, n7438, n7440, 
        \genblk1.mem_N_2584 , n7289, n7287, n7285, n7360, n7362, 
        n7364, n7366, n7368, n7370, n7372, n7374, \genblk1.mem_N_2584_adj_6030 , 
        n7294, n7296, n7298, n7300, n7302, n7304, n7306, n7308, 
        \genblk1.mem_N_2584_adj_6031 , n7217, n7215, n7339, n7337, 
        n7335;
    
    LUT4 state_2__bdd_4_lut_34641 (.A(dcache_restart_request), .B(n45183), 
         .C(state[0]), .D(state[1]), .Z(n38909)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam state_2__bdd_4_lut_34641.init = 16'ha8a0;
    FD1S3DX state_FSM_i0 (.D(n9244), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(state[2]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(476[9] 515[16])
    defparam state_FSM_i0.GSR = "ENABLED";
    FD1P3BX flush_set_i0_i0 (.D(flush_set_8__N_2513[0]), .SP(state[0]), 
            .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), .Q(flush_set[0])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam flush_set_i0_i0.GSR = "ENABLED";
    FD1P3AX refill_address__i1 (.D(\operand_m[4] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[4] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i1.GSR = "ENABLED";
    FD1S3DX refill_offset_i2 (.D(refill_offset_3__N_2489[0]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(refill_offset[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(528[5] 546[8])
    defparam refill_offset_i2.GSR = "ENABLED";
    FD1S3DX refill_request_97 (.D(refill_request_N_2565), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(dcache_refill_request)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_request_97.GSR = "ENABLED";
    FD1S3DX restart_request_99 (.D(restart_request_N_2560), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(dcache_restart_request)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam restart_request_99.GSR = "ENABLED";
    FD1S3DX refilling_93 (.D(state[2]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(dcache_refilling)) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(460[9:32])
    defparam refilling_93.GSR = "ENABLED";
    FD1S3DX state_FSM_i1 (.D(n31551), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(state[1]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(476[9] 515[16])
    defparam state_FSM_i1.GSR = "ENABLED";
    FD1S3BX state_FSM_i2 (.D(n9248), .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), 
            .Q(state[0]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(476[9] 515[16])
    defparam state_FSM_i2.GSR = "ENABLED";
    FD1P3BX flush_set_i0_i1 (.D(flush_set_8__N_2513[1]), .SP(state[0]), 
            .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), .Q(flush_set[1])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam flush_set_i0_i1.GSR = "ENABLED";
    FD1P3BX flush_set_i0_i2 (.D(flush_set_8__N_2513[2]), .SP(state[0]), 
            .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), .Q(flush_set[2])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam flush_set_i0_i2.GSR = "ENABLED";
    FD1P3BX flush_set_i0_i3 (.D(flush_set_8__N_2513[3]), .SP(state[0]), 
            .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), .Q(flush_set[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam flush_set_i0_i3.GSR = "ENABLED";
    FD1P3BX flush_set_i0_i4 (.D(flush_set_8__N_2513[4]), .SP(state[0]), 
            .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), .Q(flush_set[4])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam flush_set_i0_i4.GSR = "ENABLED";
    FD1P3BX flush_set_i0_i5 (.D(flush_set_8__N_2513[5]), .SP(state[0]), 
            .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), .Q(flush_set[5])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam flush_set_i0_i5.GSR = "ENABLED";
    FD1P3BX flush_set_i0_i6 (.D(flush_set_8__N_2513[6]), .SP(state[0]), 
            .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), .Q(flush_set[6])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam flush_set_i0_i6.GSR = "ENABLED";
    FD1P3BX flush_set_i0_i7 (.D(flush_set_8__N_2513[7]), .SP(state[0]), 
            .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), .Q(flush_set[7])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam flush_set_i0_i7.GSR = "ENABLED";
    FD1P3BX flush_set_i0_i8 (.D(flush_set_8__N_2513[8]), .SP(state[0]), 
            .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), .Q(flush_set[8])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam flush_set_i0_i8.GSR = "ENABLED";
    FD1P3AX refill_address__i2 (.D(\operand_m[5] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[5] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i2.GSR = "ENABLED";
    FD1P3AX refill_address__i3 (.D(\operand_m[6] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[6] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i3.GSR = "ENABLED";
    FD1P3AX refill_address__i4 (.D(\operand_m[7] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[7] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i4.GSR = "ENABLED";
    FD1P3AX refill_address__i5 (.D(\operand_m[8] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[8] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i5.GSR = "ENABLED";
    FD1P3AX refill_address__i6 (.D(\operand_m[9] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[9] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i6.GSR = "ENABLED";
    FD1P3AX refill_address__i7 (.D(\operand_m[10] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[10] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i7.GSR = "ENABLED";
    FD1P3AX refill_address__i8 (.D(\operand_m[11] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[11] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i8.GSR = "ENABLED";
    FD1P3AX refill_address__i9 (.D(\operand_m[12] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[12] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i9.GSR = "ENABLED";
    FD1P3AX refill_address__i10 (.D(\operand_m[13] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[13] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i10.GSR = "ENABLED";
    FD1P3AX refill_address__i11 (.D(\operand_m[14] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[14] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i11.GSR = "ENABLED";
    FD1P3AX refill_address__i12 (.D(\operand_m[15] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[15] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i12.GSR = "ENABLED";
    FD1P3AX refill_address__i13 (.D(\operand_m[16] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[16] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i13.GSR = "ENABLED";
    FD1P3AX refill_address__i14 (.D(\operand_m[17] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[17] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i14.GSR = "ENABLED";
    FD1P3AX refill_address__i15 (.D(\operand_m[18] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[18] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i15.GSR = "ENABLED";
    FD1P3AX refill_address__i16 (.D(\operand_m[19] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[19] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i16.GSR = "ENABLED";
    FD1P3AX refill_address__i17 (.D(\operand_m[20] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[20] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i17.GSR = "ENABLED";
    FD1P3AX refill_address__i18 (.D(\operand_m[21] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[21] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i18.GSR = "ENABLED";
    FD1P3AX refill_address__i19 (.D(\operand_m[22] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[22] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i19.GSR = "ENABLED";
    FD1P3AX refill_address__i20 (.D(\operand_m[23] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[23] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i20.GSR = "ENABLED";
    FD1P3AX refill_address__i21 (.D(\operand_m[24] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[24] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i21.GSR = "ENABLED";
    FD1P3AX refill_address__i22 (.D(\operand_m[25] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[25] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i22.GSR = "ENABLED";
    FD1P3AX refill_address__i23 (.D(\operand_m[26] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[26] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i23.GSR = "ENABLED";
    FD1P3AX refill_address__i24 (.D(\operand_m[27] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[27] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i24.GSR = "ENABLED";
    FD1P3AX refill_address__i25 (.D(\operand_m[28] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[28] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i25.GSR = "ENABLED";
    FD1P3AX refill_address__i26 (.D(\operand_m[29] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[29] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i26.GSR = "ENABLED";
    FD1P3AX refill_address__i27 (.D(\operand_m[30] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[30] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i27.GSR = "ENABLED";
    FD1P3AX refill_address__i28 (.D(\operand_m[31] ), .SP(REF_CLK_c_enable_1480), 
            .CK(REF_CLK_c), .Q(\dcache_refill_address[31] )) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam refill_address__i28.GSR = "ENABLED";
    FD1S3DX refill_offset_i3 (.D(refill_offset_3__N_2489[1]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(refill_offset[3])) /* synthesis LSE_LINE_FILE_ID=25, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=381, LSE_RLINE=404 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(528[5] 546[8])
    defparam refill_offset_i3.GSR = "ENABLED";
    LUT4 store_data_31__I_0_i4_3_lut (.A(store_data_m[3]), .B(wb_data_m[3]), 
         .C(state[2]), .Z(dmem_write_data[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i3_3_lut (.A(store_data_m[2]), .B(wb_data_m[2]), 
         .C(state[2]), .Z(dmem_write_data[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i5_3_lut (.A(store_data_m[4]), .B(wb_data_m[4]), 
         .C(state[2]), .Z(dmem_write_data[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(way_match_0__N_2572), .B(n45171), .C(n41284), .D(dcache_select_m), 
         .Z(miss)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(430[15:76])
    defparam i1_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_423 (.A(way_valid[0]), .B(n4), .C(n2), .D(n3), 
         .Z(way_match_0__N_2572)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(326[23:96])
    defparam i1_4_lut_adj_423.init = 16'hfffd;
    LUT4 way_tag_0__3__I_0_i4_4_lut (.A(n7540), .B(\operand_m[15] ), .C(n7541), 
         .D(n41218), .Z(n4)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A (B (C (D))+!B !(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(326[23:96])
    defparam way_tag_0__3__I_0_i4_4_lut.init = 16'h3c66;
    LUT4 way_tag_0__3__I_0_i2_4_lut (.A(n7536), .B(\operand_m[13] ), .C(n7537), 
         .D(n41218), .Z(n2)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A (B (C (D))+!B !(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(326[23:96])
    defparam way_tag_0__3__I_0_i2_4_lut.init = 16'h3c66;
    LUT4 way_tag_0__3__I_0_i3_4_lut (.A(n7538), .B(\operand_m[14] ), .C(n7539), 
         .D(n41218), .Z(n3)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A (B (C (D))+!B !(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(326[23:96])
    defparam way_tag_0__3__I_0_i3_4_lut.init = 16'h3c66;
    LUT4 store_data_31__I_0_i2_3_lut (.A(store_data_m[1]), .B(wb_data_m[1]), 
         .C(state[2]), .Z(dmem_write_data[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i1_3_lut (.A(store_data_m[0]), .B(wb_data_m[0]), 
         .C(state[2]), .Z(dmem_write_data[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 i33132_4_lut (.A(dcache_restart_request), .B(n41435), .C(icache_restart_request), 
         .D(n19852), .Z(valid_a)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+!(D))))) */ ;
    defparam i33132_4_lut.init = 16'h3233;
    LUT4 i1_4_lut_adj_424 (.A(n30107), .B(dcache_refill_ready), .C(way_match_0__N_2572), 
         .D(n41233), .Z(n9291)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(526[22:31])
    defparam i1_4_lut_adj_424.init = 16'hccce;
    LUT4 store_data_31__I_0_i24_3_lut (.A(store_data_m[23]), .B(wb_data_m[23]), 
         .C(state[2]), .Z(dmem_write_data[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i24_3_lut.init = 16'hcaca;
    LUT4 address_m_12__I_0_i1_3_lut (.A(\operand_m[2] ), .B(refill_offset[2]), 
         .C(state[2]), .Z(dmem_write_address[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(375[29] 377[63])
    defparam address_m_12__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 address_m_12__I_0_i2_3_lut (.A(\operand_m[3] ), .B(refill_offset[3]), 
         .C(state[2]), .Z(dmem_write_address[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(375[29] 377[63])
    defparam address_m_12__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 address_m_12__I_0_i3_3_lut (.A(\operand_m[4] ), .B(\dcache_refill_address[4] ), 
         .C(state[2]), .Z(dmem_write_address[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(375[29] 377[63])
    defparam address_m_12__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 address_m_12__I_0_i5_3_lut (.A(\operand_m[6] ), .B(\dcache_refill_address[6] ), 
         .C(state[2]), .Z(dmem_write_address[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(375[29] 377[63])
    defparam address_m_12__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 address_m_12__I_0_i6_3_lut (.A(\operand_m[7] ), .B(\dcache_refill_address[7] ), 
         .C(state[2]), .Z(dmem_write_address[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(375[29] 377[63])
    defparam address_m_12__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 address_m_12__I_0_i7_3_lut (.A(\operand_m[8] ), .B(\dcache_refill_address[8] ), 
         .C(state[2]), .Z(dmem_write_address[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(375[29] 377[63])
    defparam address_m_12__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 address_m_12__I_0_i10_3_lut (.A(\operand_m[11] ), .B(\dcache_refill_address[11] ), 
         .C(state[2]), .Z(dmem_write_address[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(375[29] 377[63])
    defparam address_m_12__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 address_m_12__I_0_i11_3_lut (.A(\operand_m[12] ), .B(\dcache_refill_address[12] ), 
         .C(state[2]), .Z(dmem_write_address[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(375[29] 377[63])
    defparam address_m_12__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i17_3_lut (.A(store_data_m[16]), .B(wb_data_m[16]), 
         .C(state[2]), .Z(dmem_write_data[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i17_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i18_3_lut (.A(store_data_m[17]), .B(wb_data_m[17]), 
         .C(state[2]), .Z(dmem_write_data[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i18_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i19_3_lut (.A(store_data_m[18]), .B(wb_data_m[18]), 
         .C(state[2]), .Z(dmem_write_data[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i19_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i20_3_lut (.A(store_data_m[19]), .B(wb_data_m[19]), 
         .C(state[2]), .Z(dmem_write_data[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i20_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i21_3_lut (.A(store_data_m[20]), .B(wb_data_m[20]), 
         .C(state[2]), .Z(dmem_write_data[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i21_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i22_3_lut (.A(store_data_m[21]), .B(wb_data_m[21]), 
         .C(state[2]), .Z(dmem_write_data[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i22_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i23_3_lut (.A(store_data_m[22]), .B(wb_data_m[22]), 
         .C(state[2]), .Z(dmem_write_data[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i23_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i16_3_lut (.A(store_data_m[15]), .B(wb_data_m[15]), 
         .C(state[2]), .Z(dmem_write_data[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i16_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i9_3_lut (.A(store_data_m[8]), .B(wb_data_m[8]), 
         .C(state[2]), .Z(dmem_write_data[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i10_3_lut (.A(store_data_m[9]), .B(wb_data_m[9]), 
         .C(state[2]), .Z(dmem_write_data[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i11_3_lut (.A(store_data_m[10]), .B(wb_data_m[10]), 
         .C(state[2]), .Z(dmem_write_data[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i12_3_lut (.A(store_data_m[11]), .B(wb_data_m[11]), 
         .C(state[2]), .Z(dmem_write_data[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i13_3_lut (.A(store_data_m[12]), .B(wb_data_m[12]), 
         .C(state[2]), .Z(dmem_write_data[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i13_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i14_3_lut (.A(store_data_m[13]), .B(wb_data_m[13]), 
         .C(state[2]), .Z(dmem_write_data[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i14_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i15_3_lut (.A(store_data_m[14]), .B(wb_data_m[14]), 
         .C(state[2]), .Z(dmem_write_data[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i15_3_lut.init = 16'hcaca;
    LUT4 refill_address_12__I_0_i1_3_lut (.A(\dcache_refill_address[4] ), 
         .B(flush_set[0]), .C(state[0]), .Z(tmem_write_address[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(385[29] 387[68])
    defparam refill_address_12__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 refill_address_12__I_0_i3_3_lut (.A(\dcache_refill_address[6] ), 
         .B(flush_set[2]), .C(state[0]), .Z(tmem_write_address[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(385[29] 387[68])
    defparam refill_address_12__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 refill_address_12__I_0_i4_3_lut (.A(\dcache_refill_address[7] ), 
         .B(flush_set[3]), .C(state[0]), .Z(tmem_write_address[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(385[29] 387[68])
    defparam refill_address_12__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 refill_address_12__I_0_i5_3_lut (.A(\dcache_refill_address[8] ), 
         .B(flush_set[4]), .C(state[0]), .Z(tmem_write_address[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(385[29] 387[68])
    defparam refill_address_12__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 refill_address_12__I_0_i8_3_lut (.A(\dcache_refill_address[11] ), 
         .B(flush_set[7]), .C(state[0]), .Z(tmem_write_address[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(385[29] 387[68])
    defparam refill_address_12__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 refill_address_12__I_0_i9_3_lut (.A(\dcache_refill_address[12] ), 
         .B(flush_set[8]), .C(state[0]), .Z(tmem_write_address[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(385[29] 387[68])
    defparam refill_address_12__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(state[0]), .B(dcache_refill_ready), .Z(way_tmem_we[0])) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(476[9] 515[16])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 store_data_31__I_0_i25_3_lut (.A(store_data_m[24]), .B(wb_data_m[24]), 
         .C(state[2]), .Z(dmem_write_data[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i25_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i26_3_lut (.A(store_data_m[25]), .B(wb_data_m[25]), 
         .C(state[2]), .Z(dmem_write_data[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i26_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i27_3_lut (.A(store_data_m[26]), .B(wb_data_m[26]), 
         .C(state[2]), .Z(dmem_write_data[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i27_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i28_3_lut (.A(store_data_m[27]), .B(wb_data_m[27]), 
         .C(state[2]), .Z(dmem_write_data[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i28_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i29_3_lut (.A(store_data_m[28]), .B(wb_data_m[28]), 
         .C(state[2]), .Z(dmem_write_data[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i29_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i30_3_lut (.A(store_data_m[29]), .B(wb_data_m[29]), 
         .C(state[2]), .Z(dmem_write_data[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i30_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i31_3_lut (.A(store_data_m[30]), .B(wb_data_m[30]), 
         .C(state[2]), .Z(dmem_write_data[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i31_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i32_3_lut (.A(store_data_m[31]), .B(wb_data_m[31]), 
         .C(state[2]), .Z(dmem_write_data[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i32_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_425 (.A(icache_restart_request), .B(n45183), .C(n9304), 
         .D(\state[2]_adj_181 ), .Z(n36)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(549[6:13])
    defparam i1_4_lut_adj_425.init = 16'ha8a0;
    LUT4 i1_4_lut_adj_426 (.A(n41187), .B(n41196), .C(n41203), .D(n31990), 
         .Z(n31996)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_426.init = 16'h0100;
    LUT4 i1_4_lut_adj_427 (.A(n45175), .B(way_match_0__N_2007), .C(dcache_restart_request), 
         .D(valid_f), .Z(n31990)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_427.init = 16'h0800;
    LUT4 i1_2_lut_adj_428 (.A(dcache_refill_request), .B(\operand_m[0] ), 
         .Z(\d_adr_o_31__N_2278[0] )) /* synthesis lut_function=(!(A+!(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(475[5] 516[8])
    defparam i1_2_lut_adj_428.init = 16'h4444;
    LUT4 store_data_31__I_0_i8_3_lut (.A(store_data_m[7]), .B(wb_data_m[7]), 
         .C(state[2]), .Z(dmem_write_data[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_429 (.A(state[2]), .B(refill_offset[2]), .C(dcache_refill_ready), 
         .D(n4_adj_6029), .Z(refill_offset_3__N_2489[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(529[9] 545[16])
    defparam i1_4_lut_adj_429.init = 16'hec28;
    LUT4 select_1645_Select_0_i4_4_lut (.A(dcache_refill_request), .B(state[0]), 
         .C(state[1]), .D(miss), .Z(refill_request_N_2565)) /* synthesis lut_function=(A (B+(C))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(476[9] 515[16])
    defparam select_1645_Select_0_i4_4_lut.init = 16'hf8a8;
    LUT4 i1_4_lut_adj_430 (.A(refill_offset_3__N_2557[1]), .B(refill_offset[3]), 
         .C(state[2]), .D(n4_adj_6029), .Z(refill_offset_3__N_2489[1])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(529[9] 545[16])
    defparam i1_4_lut_adj_430.init = 16'heca0;
    LUT4 i9214_3_lut (.A(refill_offset[3]), .B(refill_offset[2]), .C(dcache_refill_ready), 
         .Z(refill_offset_3__N_2557[1])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(255[5:24])
    defparam i9214_3_lut.init = 16'h6a6a;
    LUT4 i1_2_lut_rep_771 (.A(state[1]), .B(miss), .Z(n41176)) /* synthesis lut_function=(!((B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(529[9] 545[16])
    defparam i1_2_lut_rep_771.init = 16'h2222;
    LUT4 i1_3_lut_3_lut (.A(state[1]), .B(miss), .C(state[2]), .Z(n4_adj_6029)) /* synthesis lut_function=(!(A (B)+!A (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(529[9] 545[16])
    defparam i1_3_lut_3_lut.init = 16'h2727;
    LUT4 i1_3_lut_4_lut (.A(state[1]), .B(miss), .C(dflush_m), .D(n34780), 
         .Z(n31551)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(529[9] 545[16])
    defparam i1_3_lut_4_lut.init = 16'hff02;
    LUT4 i1_2_lut_rep_772 (.A(state[1]), .B(miss), .Z(REF_CLK_c_enable_1480)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(476[9] 515[16])
    defparam i1_2_lut_rep_772.init = 16'h8888;
    LUT4 i3981_3_lut_4_lut (.A(state[1]), .B(miss), .C(n41320), .D(state[2]), 
         .Z(n9244)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(476[9] 515[16])
    defparam i3981_3_lut_4_lut.init = 16'h8f88;
    LUT4 i1_4_lut_rep_773 (.A(branch_taken_m), .B(dcache_restart_request), 
         .C(n41187), .D(icache_restart_request), .Z(n41178)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(722[6:20])
    defparam i1_4_lut_rep_773.init = 16'hcdcc;
    LUT4 i33337_2_lut_4_lut (.A(branch_taken_m), .B(dcache_restart_request), 
         .C(n41187), .D(icache_restart_request), .Z(n36389)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(722[6:20])
    defparam i33337_2_lut_4_lut.init = 16'hefee;
    LUT4 i33337_rep_150_2_lut_4_lut (.A(branch_taken_m), .B(dcache_restart_request), 
         .C(n41187), .D(icache_restart_request), .Z(n37914)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(722[6:20])
    defparam i33337_rep_150_2_lut_4_lut.init = 16'hefee;
    LUT4 i33337_rep_151_2_lut_4_lut (.A(branch_taken_m), .B(dcache_restart_request), 
         .C(n41187), .D(icache_restart_request), .Z(n37915)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(722[6:20])
    defparam i33337_rep_151_2_lut_4_lut.init = 16'hefee;
    LUT4 i33337_rep_155_2_lut_4_lut (.A(branch_taken_m), .B(dcache_restart_request), 
         .C(n41187), .D(icache_restart_request), .Z(n37919)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(722[6:20])
    defparam i33337_rep_155_2_lut_4_lut.init = 16'hefee;
    LUT4 i33337_rep_153_2_lut_4_lut (.A(branch_taken_m), .B(dcache_restart_request), 
         .C(n41187), .D(icache_restart_request), .Z(n37917)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(722[6:20])
    defparam i33337_rep_153_2_lut_4_lut.init = 16'hefee;
    LUT4 i33337_rep_152_2_lut_4_lut (.A(branch_taken_m), .B(dcache_restart_request), 
         .C(n41187), .D(icache_restart_request), .Z(n37916)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(722[6:20])
    defparam i33337_rep_152_2_lut_4_lut.init = 16'hefee;
    LUT4 i33337_rep_154_2_lut_4_lut (.A(branch_taken_m), .B(dcache_restart_request), 
         .C(n41187), .D(icache_restart_request), .Z(n37918)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(722[6:20])
    defparam i33337_rep_154_2_lut_4_lut.init = 16'hefee;
    LUT4 i1_4_lut_adj_431 (.A(n23436), .B(n35822), .C(n35824), .D(n35512), 
         .Z(n34780)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(476[9] 515[16])
    defparam i1_4_lut_adj_431.init = 16'habaa;
    LUT4 i30660_4_lut (.A(flush_set[4]), .B(flush_set[6]), .C(flush_set[5]), 
         .D(flush_set[0]), .Z(n35822)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30660_4_lut.init = 16'hfffe;
    LUT4 i30662_4_lut (.A(flush_set[7]), .B(flush_set[1]), .C(flush_set[8]), 
         .D(flush_set[2]), .Z(n35824)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30662_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_432 (.A(flush_set[3]), .B(state[0]), .Z(n35512)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_432.init = 16'h4444;
    LUT4 i1_4_lut_adj_433 (.A(dflush_m), .B(state[0]), .C(n41176), .D(n31665), 
         .Z(n9248)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_433.init = 16'heca0;
    LUT4 i1_4_lut_adj_434 (.A(n35540), .B(n35538), .C(flush_set[6]), .D(flush_set[2]), 
         .Z(n31665)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_434.init = 16'hfffe;
    LUT4 i1_4_lut_adj_435 (.A(flush_set[3]), .B(flush_set[1]), .C(flush_set[8]), 
         .D(flush_set[5]), .Z(n35540)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_435.init = 16'hfffe;
    LUT4 i1_3_lut (.A(flush_set[0]), .B(flush_set[4]), .C(flush_set[7]), 
         .Z(n35538)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut.init = 16'hfefe;
    PFUMX i33552 (.BLUT(n38909), .ALUT(n38908), .C0(state[2]), .Z(restart_request_N_2560));
    LUT4 tmem_write_data_0__I_0_3_lut_4_lut (.A(refill_offset[2]), .B(refill_offset[3]), 
         .C(state[0]), .D(n30107), .Z(tmem_write_data[0])) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(193[32:45])
    defparam tmem_write_data_0__I_0_3_lut_4_lut.init = 16'h0f08;
    LUT4 state_2__bdd_2_lut_3_lut_4_lut (.A(refill_offset[2]), .B(refill_offset[3]), 
         .C(dcache_restart_request), .D(dcache_refill_ready), .Z(n38908)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(193[32:45])
    defparam state_2__bdd_2_lut_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i1_2_lut_rep_915_3_lut (.A(refill_offset[2]), .B(refill_offset[3]), 
         .C(dcache_refill_ready), .Z(n41320)) /* synthesis lut_function=(A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(193[32:45])
    defparam i1_2_lut_rep_915_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut (.A(refill_offset[2]), .B(refill_offset[3]), 
         .C(state[2]), .D(dcache_refill_ready), .Z(n23436)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(193[32:45])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    PFUMX i8 (.BLUT(n36), .ALUT(n41), .C0(icache_refill_request), .Z(restart_request_N_1998));
    LUT4 i1_2_lut_rep_767 (.A(n31996), .B(n15), .Z(n41172)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_767.init = 16'h2222;
    LUT4 i1_2_lut_3_lut (.A(n31996), .B(n15), .C(\state[2]_adj_181 ), 
         .Z(n32278)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 store_data_31__I_0_i7_3_lut (.A(store_data_m[6]), .B(wb_data_m[6]), 
         .C(state[2]), .Z(dmem_write_data[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 store_data_31__I_0_i6_3_lut (.A(store_data_m[5]), .B(wb_data_m[5]), 
         .C(state[2]), .Z(dmem_write_data[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(367[9:38])
    defparam store_data_31__I_0_i6_3_lut.init = 16'hcaca;
    \lm32_ram(data_width=32'sb0100,address_width=32'sb01001)  \memories_0..way_0_tag_ram  (.n41218(n41218), 
            .tmem_write_address({tmem_write_address[8:7], \tmem_write_address[6] , 
            \tmem_write_address[5] , tmem_write_address[4:2], \tmem_write_address[1] , 
            tmem_write_address[0]}), .n7502({n7502}), .\tmem_write_data[0] (tmem_write_data[0]), 
            .\dcache_refill_address[13] (\dcache_refill_address[13] ), .\dcache_refill_address[14] (\dcache_refill_address[14] ), 
            .\dcache_refill_address[15] (\dcache_refill_address[15] ), .n7536(n7536), 
            .n7538(n7538), .n7540(n7540), .REF_CLK_c(REF_CLK_c), .way_tmem_we({way_tmem_we}), 
            .VCC_net(VCC_net), .GND_net(GND_net), .n7541(n7541), .n7539(n7539), 
            .n7537(n7537), .\genblk1.ra ({\genblk1.ra }), .\way_valid[0] (way_valid[0])) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(299[11] 313[4])
    \lm32_ram(data_width=8,address_width=32'sb01011)  \memories_0..genblk1.byte_memories_3..way_0_data_ram  (.dmem_write_address({dmem_write_address[10:9], 
            \dmem_write_address[8] , \dmem_write_address[7] , dmem_write_address[6:4], 
            \dmem_write_address[3] , dmem_write_address[2:0]}), .n7388({n7388}), 
            .\dmem_write_data[24] (dmem_write_data[24]), .\dmem_write_data[25] (dmem_write_data[25]), 
            .\dmem_write_data[26] (dmem_write_data[26]), .\dmem_write_data[27] (dmem_write_data[27]), 
            .\dmem_write_data[28] (dmem_write_data[28]), .\dmem_write_data[29] (dmem_write_data[29]), 
            .\dmem_write_data[30] (dmem_write_data[30]), .\dmem_write_data[31] (dmem_write_data[31]), 
            .n7426(n7426), .n7428(n7428), .n7430(n7430), .n7432(n7432), 
            .n7434(n7434), .n7436(n7436), .n7438(n7438), .n7440(n7440), 
            .REF_CLK_c(REF_CLK_c), .\genblk1.mem_N_2584 (\genblk1.mem_N_2584 ), 
            .VCC_net(VCC_net), .GND_net(GND_net), .n7289(n7289), .n7287(n7287), 
            .n7285(n7285), .\byte_enable_m[3] (byte_enable_m[3]), .n9291(n9291), 
            .\state[2] (state[2]), .dcache_select_m(dcache_select_m)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(265[7] 279[7])
    \lm32_ram(data_width=8,address_width=32'sb01011)_U0  \memories_0..genblk1.byte_memories_2..way_0_data_ram  (.dmem_write_address({dmem_write_address[10:9], 
            \dmem_write_address[8] , \dmem_write_address[7] , dmem_write_address[6:4], 
            \dmem_write_address[3] , dmem_write_address[2:0]}), .n7322({n7322}), 
            .\dmem_write_data[16] (dmem_write_data[16]), .\dmem_write_data[17] (dmem_write_data[17]), 
            .\dmem_write_data[18] (dmem_write_data[18]), .\dmem_write_data[19] (dmem_write_data[19]), 
            .\dmem_write_data[20] (dmem_write_data[20]), .\dmem_write_data[21] (dmem_write_data[21]), 
            .\dmem_write_data[22] (dmem_write_data[22]), .\dmem_write_data[23] (dmem_write_data[23]), 
            .n7360(n7360), .n7362(n7362), .n7364(n7364), .n7366(n7366), 
            .n7368(n7368), .n7370(n7370), .n7372(n7372), .n7374(n7374), 
            .REF_CLK_c(REF_CLK_c), .\genblk1.mem_N_2584 (\genblk1.mem_N_2584_adj_6030 ), 
            .VCC_net(VCC_net), .GND_net(GND_net), .\byte_enable_m[2] (byte_enable_m[2]), 
            .n9291(n9291), .\state[2] (state[2]), .dcache_select_m(dcache_select_m)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(265[7] 279[7])
    \lm32_ram(data_width=8,address_width=32'sb01011)_U1  \memories_0..genblk1.byte_memories_1..way_0_data_ram  (.dmem_write_address({dmem_write_address[10:9], 
            \dmem_write_address[8] , \dmem_write_address[7] , dmem_write_address[6:4], 
            \dmem_write_address[3] , dmem_write_address[2:0]}), .n7256({n7256}), 
            .\dmem_write_data[8] (dmem_write_data[8]), .\dmem_write_data[9] (dmem_write_data[9]), 
            .\dmem_write_data[10] (dmem_write_data[10]), .\dmem_write_data[11] (dmem_write_data[11]), 
            .\dmem_write_data[12] (dmem_write_data[12]), .\dmem_write_data[13] (dmem_write_data[13]), 
            .\dmem_write_data[14] (dmem_write_data[14]), .\dmem_write_data[15] (dmem_write_data[15]), 
            .n7294(n7294), .n7296(n7296), .n7298(n7298), .n7300(n7300), 
            .n7302(n7302), .n7304(n7304), .n7306(n7306), .n7308(n7308), 
            .REF_CLK_c(REF_CLK_c), .\genblk1.mem_N_2584 (\genblk1.mem_N_2584_adj_6031 ), 
            .VCC_net(VCC_net), .GND_net(GND_net), .n7217(n7217), .n7215(n7215), 
            .n7339(n7339), .n7337(n7337), .n7335(n7335), .\byte_enable_m[1] (byte_enable_m[1]), 
            .n9291(n9291), .\state[2] (state[2]), .dcache_select_m(dcache_select_m)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(265[7] 279[7])
    \lm32_ram(data_width=8,address_width=32'sb01011)_U2  \memories_0..genblk1.byte_memories_0..way_0_data_ram  (.REF_CLK_c(REF_CLK_c), 
            .dmem_write_data({dmem_write_data}), .n7204(n7204), .n7190({n7190}), 
            .n7206(n7206), .n7208(n7208), .\genblk1.ra ({\genblk1.ra_adj_191 }), 
            .n7388({n7388}), .n7426(n7426), .n6418({n6418}), .n7224(n7224), 
            .n7289(n7289), .GND_net(GND_net), .VCC_net(VCC_net), .n7222(n7222), 
            .n7287(n7287), .n7220(n7220), .n7285(n7285), .n7428(n7428), 
            .n7430(n7430), .n7432(n7432), .n7434(n7434), .n7436(n7436), 
            .n7438(n7438), .n7440(n7440), .n7360(n7360), .n6417({n6417}), 
            .n7362(n7362), .n7364(n7364), .n7366(n7366), .\genblk1.mem_N_2584 (\genblk1.mem_N_2584_adj_6030 ), 
            .n7356(n7356), .n7322({n7322}), .n7354(n7354), .n7368(n7368), 
            .n7352(n7352), .n7350(n7350), .n7348(n7348), .n7370(n7370), 
            .n7346(n7346), .n7344(n7344), .n7342(n7342), .n7340(n7340), 
            .n7338(n7338), .n7336(n7336), .n7218(n7218), .n7372(n7372), 
            .\genblk1.mem_N_2584_adj_179 (\genblk1.mem_N_2584_adj_6031 ), 
            .n7290(n7290), .n7256({n7256}), .n7288(n7288), .n7286(n7286), 
            .n7284(n7284), .n7216(n7216), .n7374(n7374), .n7282(n7282), 
            .n7294(n7294), .n6416({n6416}), .n7296(n7296), .n7298(n7298), 
            .n7300(n7300), .n7280(n7280), .n7278(n7278), .n7214(n7214), 
            .n7302(n7302), .n7304(n7304), .n7306(n7306), .n7308(n7308), 
            .n7276(n7276), .n7274(n7274), .n7272(n7272), .dmem_write_address({dmem_write_address[10:9], 
            \dmem_write_address[8] , \dmem_write_address[7] , dmem_write_address[6:4], 
            \dmem_write_address[3] , dmem_write_address[2:0]}), .\genblk1.mem_N_2584_adj_180 (\genblk1.mem_N_2584 ), 
            .n7212(n7212), .n7270(n7270), .n7210(n7210), .n7339(n7339), 
            .n7337(n7337), .n7335(n7335), .\byte_enable_m[0] (byte_enable_m[0]), 
            .n9291(n9291), .\state[2] (state[2]), .dcache_select_m(dcache_select_m), 
            .n7217(n7217), .n7215(n7215), .dcache_data_m({dcache_data_m})) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_dcache.v(265[7] 279[7])
    
endmodule
//
// Verilog Description of module \lm32_ram(data_width=32'sb0100,address_width=32'sb01001) 
//

module \lm32_ram(data_width=32'sb0100,address_width=32'sb01001)  (n41218, 
            tmem_write_address, n7502, \tmem_write_data[0] , \dcache_refill_address[13] , 
            \dcache_refill_address[14] , \dcache_refill_address[15] , n7536, 
            n7538, n7540, REF_CLK_c, way_tmem_we, VCC_net, GND_net, 
            n7541, n7539, n7537, \genblk1.ra , \way_valid[0] ) /* synthesis syn_module_defined=1 */ ;
    output n41218;
    input [8:0]tmem_write_address;
    input [8:0]n7502;
    input \tmem_write_data[0] ;
    input \dcache_refill_address[13] ;
    input \dcache_refill_address[14] ;
    input \dcache_refill_address[15] ;
    output n7536;
    output n7538;
    output n7540;
    input REF_CLK_c;
    input [0:0]way_tmem_we;
    input VCC_net;
    input GND_net;
    output n7541;
    output n7539;
    output n7537;
    output [8:0]\genblk1.ra ;
    output \way_valid[0] ;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    
    wire n7532, n7531, n7534, n7535, n7529, n7527, n7525, n7523, 
        n7521, n7519, n7517, n7515, n7513, n27373, n27372;
    
    LUT4 i3136_2_lut_rep_813 (.A(n7532), .B(n7531), .Z(n41218)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam i3136_2_lut_rep_813.init = 16'h8888;
    DP16KD \genblk1.mem0  (.DIA0(\tmem_write_data[0] ), .DIA1(\dcache_refill_address[13] ), 
           .DIA2(\dcache_refill_address[14] ), .DIA3(\dcache_refill_address[15] ), 
           .DIA4(GND_net), .DIA5(GND_net), .DIA6(GND_net), .DIA7(GND_net), 
           .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), .DIA11(GND_net), 
           .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), .DIA15(GND_net), 
           .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), .ADA1(GND_net), 
           .ADA2(tmem_write_address[0]), .ADA3(tmem_write_address[1]), .ADA4(tmem_write_address[2]), 
           .ADA5(tmem_write_address[3]), .ADA6(tmem_write_address[4]), .ADA7(tmem_write_address[5]), 
           .ADA8(tmem_write_address[6]), .ADA9(tmem_write_address[7]), .ADA10(tmem_write_address[8]), 
           .ADA11(GND_net), .ADA12(GND_net), .ADA13(GND_net), .CEA(VCC_net), 
           .OCEA(VCC_net), .CLKA(REF_CLK_c), .WEA(way_tmem_we[0]), .CSA0(GND_net), 
           .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), 
           .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
           .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
           .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), .DIB12(GND_net), 
           .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), .DIB16(GND_net), 
           .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(n7502[0]), 
           .ADB3(n7502[1]), .ADB4(n7502[2]), .ADB5(n7502[3]), .ADB6(n7502[4]), 
           .ADB7(n7502[5]), .ADB8(n7502[6]), .ADB9(n7502[7]), .ADB10(n7502[8]), 
           .ADB11(GND_net), .ADB12(GND_net), .ADB13(GND_net), .CEB(VCC_net), 
           .OCEB(VCC_net), .CLKB(REF_CLK_c), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(GND_net), .DOB0(n7534), 
           .DOB1(n7536), .DOB2(n7538), .DOB3(n7540));
    defparam \genblk1.mem0 .DATA_WIDTH_A = 4;
    defparam \genblk1.mem0 .DATA_WIDTH_B = 4;
    defparam \genblk1.mem0 .REGMODE_A = "NOREG";
    defparam \genblk1.mem0 .REGMODE_B = "NOREG";
    defparam \genblk1.mem0 .RESETMODE = "SYNC";
    defparam \genblk1.mem0 .ASYNC_RESET_RELEASE = "SYNC";
    defparam \genblk1.mem0 .WRITEMODE_A = "WRITETHROUGH";
    defparam \genblk1.mem0 .WRITEMODE_B = "WRITETHROUGH";
    defparam \genblk1.mem0 .CSDECODE_A = "0b000";
    defparam \genblk1.mem0 .CSDECODE_B = "0b000";
    defparam \genblk1.mem0 .GSR = "DISABLED";
    defparam \genblk1.mem0 .INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INIT_DATA = "STATIC";
    FD1S3AX \genblk1.mem  (.D(\dcache_refill_address[15] ), .CK(REF_CLK_c), 
            .Q(n7541));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3140  (.D(\dcache_refill_address[14] ), .CK(REF_CLK_c), 
            .Q(n7539));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3140 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3139  (.D(\dcache_refill_address[13] ), .CK(REF_CLK_c), 
            .Q(n7537));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3139 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3138  (.D(\tmem_write_data[0] ), .CK(REF_CLK_c), 
            .Q(n7535));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3138 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3137  (.D(way_tmem_we[0]), .CK(REF_CLK_c), .Q(n7532));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3137 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3135  (.D(n7502[8]), .CK(REF_CLK_c), .Q(\genblk1.ra [8]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3135 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3133  (.D(tmem_write_address[8]), .CK(REF_CLK_c), 
            .Q(n7529));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3133 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3132  (.D(n7502[7]), .CK(REF_CLK_c), .Q(\genblk1.ra [7]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3132 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3131  (.D(tmem_write_address[7]), .CK(REF_CLK_c), 
            .Q(n7527));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3131 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3130  (.D(n7502[6]), .CK(REF_CLK_c), .Q(\genblk1.ra [6]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3130 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3129  (.D(tmem_write_address[6]), .CK(REF_CLK_c), 
            .Q(n7525));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3129 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3128  (.D(n7502[5]), .CK(REF_CLK_c), .Q(\genblk1.ra [5]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3128 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3127  (.D(tmem_write_address[5]), .CK(REF_CLK_c), 
            .Q(n7523));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3127 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3126  (.D(n7502[4]), .CK(REF_CLK_c), .Q(\genblk1.ra [4]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3126 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3125  (.D(tmem_write_address[4]), .CK(REF_CLK_c), 
            .Q(n7521));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3125 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3124  (.D(n7502[3]), .CK(REF_CLK_c), .Q(\genblk1.ra [3]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3124 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3123  (.D(tmem_write_address[3]), .CK(REF_CLK_c), 
            .Q(n7519));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3123 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3122  (.D(n7502[2]), .CK(REF_CLK_c), .Q(\genblk1.ra [2]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3122 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3121  (.D(tmem_write_address[2]), .CK(REF_CLK_c), 
            .Q(n7517));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3121 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3120  (.D(n7502[1]), .CK(REF_CLK_c), .Q(\genblk1.ra [1]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3120 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3119  (.D(tmem_write_address[1]), .CK(REF_CLK_c), 
            .Q(n7515));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3119 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3118  (.D(n7502[0]), .CK(REF_CLK_c), .Q(\genblk1.ra [0]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3118 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3117  (.D(tmem_write_address[0]), .CK(REF_CLK_c), 
            .Q(n7513));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3117 .GSR = "ENABLED";
    LUT4 mux_3140_i1_3_lut_4_lut (.A(n7532), .B(n7531), .C(n7535), .D(n7534), 
         .Z(\way_valid[0] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3140_i1_3_lut_4_lut.init = 16'hf780;
    CCU2C equal_3133_9 (.A0(\genblk1.ra [1]), .B0(n7515), .C0(\genblk1.ra [0]), 
          .D0(n7513), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27373), .S1(n7531));
    defparam equal_3133_9.INIT0 = 16'h9009;
    defparam equal_3133_9.INIT1 = 16'h0000;
    defparam equal_3133_9.INJECT1_0 = "YES";
    defparam equal_3133_9.INJECT1_1 = "NO";
    CCU2C equal_3133_8 (.A0(\genblk1.ra [5]), .B0(n7523), .C0(\genblk1.ra [4]), 
          .D0(n7521), .A1(\genblk1.ra [3]), .B1(n7519), .C1(\genblk1.ra [2]), 
          .D1(n7517), .CIN(n27372), .COUT(n27373));
    defparam equal_3133_8.INIT0 = 16'h9009;
    defparam equal_3133_8.INIT1 = 16'h9009;
    defparam equal_3133_8.INJECT1_0 = "YES";
    defparam equal_3133_8.INJECT1_1 = "YES";
    CCU2C equal_3133_0 (.A0(\genblk1.ra [8]), .B0(n7529), .C0(GND_net), 
          .D0(VCC_net), .A1(\genblk1.ra [7]), .B1(n7527), .C1(\genblk1.ra [6]), 
          .D1(n7525), .COUT(n27372));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam equal_3133_0.INIT0 = 16'h0009;
    defparam equal_3133_0.INIT1 = 16'h9009;
    defparam equal_3133_0.INJECT1_0 = "NO";
    defparam equal_3133_0.INJECT1_1 = "YES";
    
endmodule
//
// Verilog Description of module \lm32_ram(data_width=8,address_width=32'sb01011) 
//

module \lm32_ram(data_width=8,address_width=32'sb01011)  (dmem_write_address, 
            n7388, \dmem_write_data[24] , \dmem_write_data[25] , \dmem_write_data[26] , 
            \dmem_write_data[27] , \dmem_write_data[28] , \dmem_write_data[29] , 
            \dmem_write_data[30] , \dmem_write_data[31] , n7426, n7428, 
            n7430, n7432, n7434, n7436, n7438, n7440, REF_CLK_c, 
            \genblk1.mem_N_2584 , VCC_net, GND_net, n7289, n7287, 
            n7285, \byte_enable_m[3] , n9291, \state[2] , dcache_select_m) /* synthesis syn_module_defined=1 */ ;
    input [10:0]dmem_write_address;
    input [10:0]n7388;
    input \dmem_write_data[24] ;
    input \dmem_write_data[25] ;
    input \dmem_write_data[26] ;
    input \dmem_write_data[27] ;
    input \dmem_write_data[28] ;
    input \dmem_write_data[29] ;
    input \dmem_write_data[30] ;
    input \dmem_write_data[31] ;
    output n7426;
    output n7428;
    output n7430;
    output n7432;
    output n7434;
    output n7436;
    output n7438;
    output n7440;
    input REF_CLK_c;
    output \genblk1.mem_N_2584 ;
    input VCC_net;
    input GND_net;
    output n7289;
    output n7287;
    output n7285;
    input \byte_enable_m[3] ;
    input n9291;
    input \state[2] ;
    input dcache_select_m;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    
    DP16KD \genblk1.mem0  (.DIA0(\dmem_write_data[24] ), .DIA1(\dmem_write_data[25] ), 
           .DIA2(\dmem_write_data[26] ), .DIA3(\dmem_write_data[27] ), .DIA4(\dmem_write_data[28] ), 
           .DIA5(\dmem_write_data[29] ), .DIA6(\dmem_write_data[30] ), .DIA7(\dmem_write_data[31] ), 
           .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), .DIA11(GND_net), 
           .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), .DIA15(GND_net), 
           .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), .ADA1(GND_net), 
           .ADA2(GND_net), .ADA3(dmem_write_address[0]), .ADA4(dmem_write_address[1]), 
           .ADA5(dmem_write_address[2]), .ADA6(dmem_write_address[3]), .ADA7(dmem_write_address[4]), 
           .ADA8(dmem_write_address[5]), .ADA9(dmem_write_address[6]), .ADA10(dmem_write_address[7]), 
           .ADA11(dmem_write_address[8]), .ADA12(dmem_write_address[9]), 
           .ADA13(dmem_write_address[10]), .CEA(VCC_net), .OCEA(VCC_net), 
           .CLKA(REF_CLK_c), .WEA(\genblk1.mem_N_2584 ), .CSA0(GND_net), 
           .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), 
           .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
           .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
           .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), .DIB12(GND_net), 
           .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), .DIB16(GND_net), 
           .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
           .ADB3(n7388[0]), .ADB4(n7388[1]), .ADB5(n7388[2]), .ADB6(n7388[3]), 
           .ADB7(n7388[4]), .ADB8(n7388[5]), .ADB9(n7388[6]), .ADB10(n7388[7]), 
           .ADB11(n7388[8]), .ADB12(n7388[9]), .ADB13(n7388[10]), .CEB(VCC_net), 
           .OCEB(VCC_net), .CLKB(REF_CLK_c), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(GND_net), .DOB0(n7426), 
           .DOB1(n7428), .DOB2(n7430), .DOB3(n7432), .DOB4(n7434), .DOB5(n7436), 
           .DOB6(n7438), .DOB7(n7440));
    defparam \genblk1.mem0 .DATA_WIDTH_A = 9;
    defparam \genblk1.mem0 .DATA_WIDTH_B = 9;
    defparam \genblk1.mem0 .REGMODE_A = "NOREG";
    defparam \genblk1.mem0 .REGMODE_B = "NOREG";
    defparam \genblk1.mem0 .RESETMODE = "SYNC";
    defparam \genblk1.mem0 .ASYNC_RESET_RELEASE = "SYNC";
    defparam \genblk1.mem0 .WRITEMODE_A = "WRITETHROUGH";
    defparam \genblk1.mem0 .WRITEMODE_B = "WRITETHROUGH";
    defparam \genblk1.mem0 .CSDECODE_A = "0b000";
    defparam \genblk1.mem0 .CSDECODE_B = "0b000";
    defparam \genblk1.mem0 .GSR = "DISABLED";
    defparam \genblk1.mem0 .INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INIT_DATA = "STATIC";
    FD1S3AX \genblk1.mem_3077  (.D(dmem_write_address[10]), .CK(REF_CLK_c), 
            .Q(n7289));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3077 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3075  (.D(dmem_write_address[9]), .CK(REF_CLK_c), 
            .Q(n7287));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3075 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3073  (.D(dmem_write_address[8]), .CK(REF_CLK_c), 
            .Q(n7285));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3073 .GSR = "ENABLED";
    LUT4 i2_4_lut (.A(\byte_enable_m[3] ), .B(n9291), .C(\state[2] ), 
         .D(dcache_select_m), .Z(\genblk1.mem_N_2584 )) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(298[13:63])
    defparam i2_4_lut.init = 16'hc8c0;
    
endmodule
//
// Verilog Description of module \lm32_ram(data_width=8,address_width=32'sb01011)_U0 
//

module \lm32_ram(data_width=8,address_width=32'sb01011)_U0  (dmem_write_address, 
            n7322, \dmem_write_data[16] , \dmem_write_data[17] , \dmem_write_data[18] , 
            \dmem_write_data[19] , \dmem_write_data[20] , \dmem_write_data[21] , 
            \dmem_write_data[22] , \dmem_write_data[23] , n7360, n7362, 
            n7364, n7366, n7368, n7370, n7372, n7374, REF_CLK_c, 
            \genblk1.mem_N_2584 , VCC_net, GND_net, \byte_enable_m[2] , 
            n9291, \state[2] , dcache_select_m) /* synthesis syn_module_defined=1 */ ;
    input [10:0]dmem_write_address;
    input [10:0]n7322;
    input \dmem_write_data[16] ;
    input \dmem_write_data[17] ;
    input \dmem_write_data[18] ;
    input \dmem_write_data[19] ;
    input \dmem_write_data[20] ;
    input \dmem_write_data[21] ;
    input \dmem_write_data[22] ;
    input \dmem_write_data[23] ;
    output n7360;
    output n7362;
    output n7364;
    output n7366;
    output n7368;
    output n7370;
    output n7372;
    output n7374;
    input REF_CLK_c;
    output \genblk1.mem_N_2584 ;
    input VCC_net;
    input GND_net;
    input \byte_enable_m[2] ;
    input n9291;
    input \state[2] ;
    input dcache_select_m;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    
    DP16KD \genblk1.mem0  (.DIA0(\dmem_write_data[16] ), .DIA1(\dmem_write_data[17] ), 
           .DIA2(\dmem_write_data[18] ), .DIA3(\dmem_write_data[19] ), .DIA4(\dmem_write_data[20] ), 
           .DIA5(\dmem_write_data[21] ), .DIA6(\dmem_write_data[22] ), .DIA7(\dmem_write_data[23] ), 
           .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), .DIA11(GND_net), 
           .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), .DIA15(GND_net), 
           .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), .ADA1(GND_net), 
           .ADA2(GND_net), .ADA3(dmem_write_address[0]), .ADA4(dmem_write_address[1]), 
           .ADA5(dmem_write_address[2]), .ADA6(dmem_write_address[3]), .ADA7(dmem_write_address[4]), 
           .ADA8(dmem_write_address[5]), .ADA9(dmem_write_address[6]), .ADA10(dmem_write_address[7]), 
           .ADA11(dmem_write_address[8]), .ADA12(dmem_write_address[9]), 
           .ADA13(dmem_write_address[10]), .CEA(VCC_net), .OCEA(VCC_net), 
           .CLKA(REF_CLK_c), .WEA(\genblk1.mem_N_2584 ), .CSA0(GND_net), 
           .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), 
           .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
           .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
           .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), .DIB12(GND_net), 
           .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), .DIB16(GND_net), 
           .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
           .ADB3(n7322[0]), .ADB4(n7322[1]), .ADB5(n7322[2]), .ADB6(n7322[3]), 
           .ADB7(n7322[4]), .ADB8(n7322[5]), .ADB9(n7322[6]), .ADB10(n7322[7]), 
           .ADB11(n7322[8]), .ADB12(n7322[9]), .ADB13(n7322[10]), .CEB(VCC_net), 
           .OCEB(VCC_net), .CLKB(REF_CLK_c), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(GND_net), .DOB0(n7360), 
           .DOB1(n7362), .DOB2(n7364), .DOB3(n7366), .DOB4(n7368), .DOB5(n7370), 
           .DOB6(n7372), .DOB7(n7374));
    defparam \genblk1.mem0 .DATA_WIDTH_A = 9;
    defparam \genblk1.mem0 .DATA_WIDTH_B = 9;
    defparam \genblk1.mem0 .REGMODE_A = "NOREG";
    defparam \genblk1.mem0 .REGMODE_B = "NOREG";
    defparam \genblk1.mem0 .RESETMODE = "SYNC";
    defparam \genblk1.mem0 .ASYNC_RESET_RELEASE = "SYNC";
    defparam \genblk1.mem0 .WRITEMODE_A = "WRITETHROUGH";
    defparam \genblk1.mem0 .WRITEMODE_B = "WRITETHROUGH";
    defparam \genblk1.mem0 .CSDECODE_A = "0b000";
    defparam \genblk1.mem0 .CSDECODE_B = "0b000";
    defparam \genblk1.mem0 .GSR = "DISABLED";
    defparam \genblk1.mem0 .INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INIT_DATA = "STATIC";
    LUT4 i2_4_lut (.A(\byte_enable_m[2] ), .B(n9291), .C(\state[2] ), 
         .D(dcache_select_m), .Z(\genblk1.mem_N_2584 )) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(298[13:63])
    defparam i2_4_lut.init = 16'hc8c0;
    
endmodule
//
// Verilog Description of module \lm32_ram(data_width=8,address_width=32'sb01011)_U1 
//

module \lm32_ram(data_width=8,address_width=32'sb01011)_U1  (dmem_write_address, 
            n7256, \dmem_write_data[8] , \dmem_write_data[9] , \dmem_write_data[10] , 
            \dmem_write_data[11] , \dmem_write_data[12] , \dmem_write_data[13] , 
            \dmem_write_data[14] , \dmem_write_data[15] , n7294, n7296, 
            n7298, n7300, n7302, n7304, n7306, n7308, REF_CLK_c, 
            \genblk1.mem_N_2584 , VCC_net, GND_net, n7217, n7215, 
            n7339, n7337, n7335, \byte_enable_m[1] , n9291, \state[2] , 
            dcache_select_m) /* synthesis syn_module_defined=1 */ ;
    input [10:0]dmem_write_address;
    input [10:0]n7256;
    input \dmem_write_data[8] ;
    input \dmem_write_data[9] ;
    input \dmem_write_data[10] ;
    input \dmem_write_data[11] ;
    input \dmem_write_data[12] ;
    input \dmem_write_data[13] ;
    input \dmem_write_data[14] ;
    input \dmem_write_data[15] ;
    output n7294;
    output n7296;
    output n7298;
    output n7300;
    output n7302;
    output n7304;
    output n7306;
    output n7308;
    input REF_CLK_c;
    output \genblk1.mem_N_2584 ;
    input VCC_net;
    input GND_net;
    output n7217;
    output n7215;
    output n7339;
    output n7337;
    output n7335;
    input \byte_enable_m[1] ;
    input n9291;
    input \state[2] ;
    input dcache_select_m;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    
    DP16KD \genblk1.mem0  (.DIA0(\dmem_write_data[8] ), .DIA1(\dmem_write_data[9] ), 
           .DIA2(\dmem_write_data[10] ), .DIA3(\dmem_write_data[11] ), .DIA4(\dmem_write_data[12] ), 
           .DIA5(\dmem_write_data[13] ), .DIA6(\dmem_write_data[14] ), .DIA7(\dmem_write_data[15] ), 
           .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), .DIA11(GND_net), 
           .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), .DIA15(GND_net), 
           .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), .ADA1(GND_net), 
           .ADA2(GND_net), .ADA3(dmem_write_address[0]), .ADA4(dmem_write_address[1]), 
           .ADA5(dmem_write_address[2]), .ADA6(dmem_write_address[3]), .ADA7(dmem_write_address[4]), 
           .ADA8(dmem_write_address[5]), .ADA9(dmem_write_address[6]), .ADA10(dmem_write_address[7]), 
           .ADA11(dmem_write_address[8]), .ADA12(dmem_write_address[9]), 
           .ADA13(dmem_write_address[10]), .CEA(VCC_net), .OCEA(VCC_net), 
           .CLKA(REF_CLK_c), .WEA(\genblk1.mem_N_2584 ), .CSA0(GND_net), 
           .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), 
           .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
           .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
           .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), .DIB12(GND_net), 
           .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), .DIB16(GND_net), 
           .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
           .ADB3(n7256[0]), .ADB4(n7256[1]), .ADB5(n7256[2]), .ADB6(n7256[3]), 
           .ADB7(n7256[4]), .ADB8(n7256[5]), .ADB9(n7256[6]), .ADB10(n7256[7]), 
           .ADB11(n7256[8]), .ADB12(n7256[9]), .ADB13(n7256[10]), .CEB(VCC_net), 
           .OCEB(VCC_net), .CLKB(REF_CLK_c), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(GND_net), .DOB0(n7294), 
           .DOB1(n7296), .DOB2(n7298), .DOB3(n7300), .DOB4(n7302), .DOB5(n7304), 
           .DOB6(n7306), .DOB7(n7308));
    defparam \genblk1.mem0 .DATA_WIDTH_A = 9;
    defparam \genblk1.mem0 .DATA_WIDTH_B = 9;
    defparam \genblk1.mem0 .REGMODE_A = "NOREG";
    defparam \genblk1.mem0 .REGMODE_B = "NOREG";
    defparam \genblk1.mem0 .RESETMODE = "SYNC";
    defparam \genblk1.mem0 .ASYNC_RESET_RELEASE = "SYNC";
    defparam \genblk1.mem0 .WRITEMODE_A = "WRITETHROUGH";
    defparam \genblk1.mem0 .WRITEMODE_B = "WRITETHROUGH";
    defparam \genblk1.mem0 .CSDECODE_A = "0b000";
    defparam \genblk1.mem0 .CSDECODE_B = "0b000";
    defparam \genblk1.mem0 .GSR = "DISABLED";
    defparam \genblk1.mem0 .INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INIT_DATA = "STATIC";
    FD1S3AX \genblk1.mem_3003  (.D(dmem_write_address[7]), .CK(REF_CLK_c), 
            .Q(n7217));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3003 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3001  (.D(dmem_write_address[6]), .CK(REF_CLK_c), 
            .Q(n7215));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3001 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2993  (.D(dmem_write_address[2]), .CK(REF_CLK_c), 
            .Q(n7339));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_2993 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2991  (.D(dmem_write_address[1]), .CK(REF_CLK_c), 
            .Q(n7337));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_2991 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2989  (.D(dmem_write_address[0]), .CK(REF_CLK_c), 
            .Q(n7335));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_2989 .GSR = "ENABLED";
    LUT4 i2_4_lut (.A(\byte_enable_m[1] ), .B(n9291), .C(\state[2] ), 
         .D(dcache_select_m), .Z(\genblk1.mem_N_2584 )) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(298[13:63])
    defparam i2_4_lut.init = 16'hc8c0;
    
endmodule
//
// Verilog Description of module \lm32_ram(data_width=8,address_width=32'sb01011)_U2 
//

module \lm32_ram(data_width=8,address_width=32'sb01011)_U2  (REF_CLK_c, dmem_write_data, 
            n7204, n7190, n7206, n7208, \genblk1.ra , n7388, n7426, 
            n6418, n7224, n7289, GND_net, VCC_net, n7222, n7287, 
            n7220, n7285, n7428, n7430, n7432, n7434, n7436, n7438, 
            n7440, n7360, n6417, n7362, n7364, n7366, \genblk1.mem_N_2584 , 
            n7356, n7322, n7354, n7368, n7352, n7350, n7348, n7370, 
            n7346, n7344, n7342, n7340, n7338, n7336, n7218, n7372, 
            \genblk1.mem_N_2584_adj_179 , n7290, n7256, n7288, n7286, 
            n7284, n7216, n7374, n7282, n7294, n6416, n7296, n7298, 
            n7300, n7280, n7278, n7214, n7302, n7304, n7306, n7308, 
            n7276, n7274, n7272, dmem_write_address, \genblk1.mem_N_2584_adj_180 , 
            n7212, n7270, n7210, n7339, n7337, n7335, \byte_enable_m[0] , 
            n9291, \state[2] , dcache_select_m, n7217, n7215, dcache_data_m) /* synthesis syn_module_defined=1 */ ;
    input REF_CLK_c;
    input [31:0]dmem_write_data;
    output n7204;
    input [10:0]n7190;
    output n7206;
    output n7208;
    output [10:0]\genblk1.ra ;
    input [10:0]n7388;
    input n7426;
    output [7:0]n6418;
    output n7224;
    input n7289;
    input GND_net;
    input VCC_net;
    output n7222;
    input n7287;
    output n7220;
    input n7285;
    input n7428;
    input n7430;
    input n7432;
    input n7434;
    input n7436;
    input n7438;
    input n7440;
    input n7360;
    output [7:0]n6417;
    input n7362;
    input n7364;
    input n7366;
    input \genblk1.mem_N_2584 ;
    output n7356;
    input [10:0]n7322;
    output n7354;
    input n7368;
    output n7352;
    output n7350;
    output n7348;
    input n7370;
    output n7346;
    output n7344;
    output n7342;
    output n7340;
    output n7338;
    output n7336;
    output n7218;
    input n7372;
    input \genblk1.mem_N_2584_adj_179 ;
    output n7290;
    input [10:0]n7256;
    output n7288;
    output n7286;
    output n7284;
    output n7216;
    input n7374;
    output n7282;
    input n7294;
    output [7:0]n6416;
    input n7296;
    input n7298;
    input n7300;
    output n7280;
    output n7278;
    output n7214;
    input n7302;
    input n7304;
    input n7306;
    input n7308;
    output n7276;
    output n7274;
    output n7272;
    input [10:0]dmem_write_address;
    input \genblk1.mem_N_2584_adj_180 ;
    output n7212;
    output n7270;
    output n7210;
    input n7339;
    input n7337;
    input n7335;
    input \byte_enable_m[0] ;
    input n9291;
    input \state[2] ;
    input dcache_select_m;
    input n7217;
    input n7215;
    output [7:0]dcache_data_m;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    
    wire n7241, n7239, n7237, n7235, n7233, n7231, n7229, n7424, 
        n7423, n7427, n27366, n7429, n7431, n7433, n7435, n7437, 
        n7439, n7441, n7358, n7357, n7361, n7363, n7365, n7367, 
        n7226, \genblk1.mem_N_2584_c , n7375, n7373, n7371, n7369, 
        n7309, n7307, n7305, n7303, n7301, n7299, n7297, n7295, 
        n7292, n7291, n7279, n7277, n7228, n7230, n7232, n7234, 
        n7236, n7238, n7240, n7242, n7243, n27381, n7275, n27380, 
        n27379, n27378, n27377, n27376, n7225, n27371, n27370, 
        n27369, n27368, n27367;
    
    FD1S3AX \genblk1.mem_2986  (.D(dmem_write_data[6]), .CK(REF_CLK_c), 
            .Q(n7241));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2986 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2985  (.D(dmem_write_data[5]), .CK(REF_CLK_c), 
            .Q(n7239));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2985 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2984  (.D(dmem_write_data[4]), .CK(REF_CLK_c), 
            .Q(n7237));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2984 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2956  (.D(n7190[0]), .CK(REF_CLK_c), .Q(n7204));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2956 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2958  (.D(n7190[1]), .CK(REF_CLK_c), .Q(n7206));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2958 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2960  (.D(n7190[2]), .CK(REF_CLK_c), .Q(n7208));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2960 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2983  (.D(dmem_write_data[3]), .CK(REF_CLK_c), 
            .Q(n7235));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2983 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2982  (.D(dmem_write_data[2]), .CK(REF_CLK_c), 
            .Q(n7233));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2982 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3070  (.D(n7388[6]), .CK(REF_CLK_c), .Q(\genblk1.ra [6]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3070 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3068  (.D(n7388[5]), .CK(REF_CLK_c), .Q(\genblk1.ra [5]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3068 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3066  (.D(n7388[4]), .CK(REF_CLK_c), .Q(\genblk1.ra [4]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3066 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3064  (.D(n7388[3]), .CK(REF_CLK_c), .Q(\genblk1.ra [3]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3064 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2981  (.D(dmem_write_data[1]), .CK(REF_CLK_c), 
            .Q(n7231));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2981 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2980  (.D(dmem_write_data[0]), .CK(REF_CLK_c), 
            .Q(n7229));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2980 .GSR = "ENABLED";
    LUT4 mux_3088_i1_3_lut_4_lut (.A(n7424), .B(n7423), .C(n7427), .D(n7426), 
         .Z(n6418[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3088_i1_3_lut_4_lut.init = 16'hf780;
    CCU2C equal_2975_0 (.A0(n7224), .B0(n7289), .C0(GND_net), .D0(VCC_net), 
          .A1(n7222), .B1(n7287), .C1(n7220), .D1(n7285), .COUT(n27366));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam equal_2975_0.INIT0 = 16'h0009;
    defparam equal_2975_0.INIT1 = 16'h9009;
    defparam equal_2975_0.INJECT1_0 = "NO";
    defparam equal_2975_0.INJECT1_1 = "YES";
    FD1S3AX \genblk1.mem_3062  (.D(n7388[2]), .CK(REF_CLK_c), .Q(\genblk1.ra [2]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3062 .GSR = "ENABLED";
    LUT4 mux_3088_i2_3_lut_4_lut (.A(n7424), .B(n7423), .C(n7429), .D(n7428), 
         .Z(n6418[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3088_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3088_i3_3_lut_4_lut (.A(n7424), .B(n7423), .C(n7431), .D(n7430), 
         .Z(n6418[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3088_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3088_i4_3_lut_4_lut (.A(n7424), .B(n7423), .C(n7433), .D(n7432), 
         .Z(n6418[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3088_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3088_i5_3_lut_4_lut (.A(n7424), .B(n7423), .C(n7435), .D(n7434), 
         .Z(n6418[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3088_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3088_i6_3_lut_4_lut (.A(n7424), .B(n7423), .C(n7437), .D(n7436), 
         .Z(n6418[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3088_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3088_i7_3_lut_4_lut (.A(n7424), .B(n7423), .C(n7439), .D(n7438), 
         .Z(n6418[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3088_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3088_i8_3_lut_4_lut (.A(n7424), .B(n7423), .C(n7441), .D(n7440), 
         .Z(n6418[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3088_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3054_i1_3_lut_4_lut (.A(n7358), .B(n7357), .C(n7361), .D(n7360), 
         .Z(n6417[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3054_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3054_i2_3_lut_4_lut (.A(n7358), .B(n7357), .C(n7363), .D(n7362), 
         .Z(n6417[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3054_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3054_i3_3_lut_4_lut (.A(n7358), .B(n7357), .C(n7365), .D(n7364), 
         .Z(n6417[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3054_i3_3_lut_4_lut.init = 16'hf780;
    FD1S3AX \genblk1.mem_3060  (.D(n7388[1]), .CK(REF_CLK_c), .Q(\genblk1.ra [1]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3060 .GSR = "ENABLED";
    LUT4 mux_3054_i4_3_lut_4_lut (.A(n7358), .B(n7357), .C(n7367), .D(n7366), 
         .Z(n6417[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3054_i4_3_lut_4_lut.init = 16'hf780;
    FD1S3AX \genblk1.mem_2979  (.D(\genblk1.mem_N_2584_c ), .CK(REF_CLK_c), 
            .Q(n7226));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2979 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2977  (.D(n7190[10]), .CK(REF_CLK_c), .Q(n7224));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2977 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2974  (.D(n7190[9]), .CK(REF_CLK_c), .Q(n7222));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2974 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3058  (.D(n7388[0]), .CK(REF_CLK_c), .Q(\genblk1.ra [0]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3058 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem  (.D(dmem_write_data[23]), .CK(REF_CLK_c), .Q(n7375));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3054  (.D(dmem_write_data[22]), .CK(REF_CLK_c), 
            .Q(n7373));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3054 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3053  (.D(dmem_write_data[21]), .CK(REF_CLK_c), 
            .Q(n7371));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3053 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3052  (.D(dmem_write_data[20]), .CK(REF_CLK_c), 
            .Q(n7369));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3052 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3051  (.D(dmem_write_data[19]), .CK(REF_CLK_c), 
            .Q(n7367));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3051 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3050  (.D(dmem_write_data[18]), .CK(REF_CLK_c), 
            .Q(n7365));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3050 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3049  (.D(dmem_write_data[17]), .CK(REF_CLK_c), 
            .Q(n7363));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3049 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3048  (.D(dmem_write_data[16]), .CK(REF_CLK_c), 
            .Q(n7361));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3048 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3047  (.D(\genblk1.mem_N_2584 ), .CK(REF_CLK_c), 
            .Q(n7358));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3047 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3045  (.D(n7322[10]), .CK(REF_CLK_c), .Q(n7356));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3045 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3042  (.D(n7322[9]), .CK(REF_CLK_c), .Q(n7354));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3042 .GSR = "ENABLED";
    LUT4 mux_3054_i5_3_lut_4_lut (.A(n7358), .B(n7357), .C(n7369), .D(n7368), 
         .Z(n6417[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3054_i5_3_lut_4_lut.init = 16'hf780;
    FD1S3AX \genblk1.mem_3040  (.D(n7322[8]), .CK(REF_CLK_c), .Q(n7352));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3040 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3038  (.D(n7322[7]), .CK(REF_CLK_c), .Q(n7350));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3038 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3036  (.D(n7322[6]), .CK(REF_CLK_c), .Q(n7348));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3036 .GSR = "ENABLED";
    LUT4 mux_3054_i6_3_lut_4_lut (.A(n7358), .B(n7357), .C(n7371), .D(n7370), 
         .Z(n6417[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3054_i6_3_lut_4_lut.init = 16'hf780;
    FD1S3AX \genblk1.mem_3034  (.D(n7322[5]), .CK(REF_CLK_c), .Q(n7346));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3034 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3032  (.D(n7322[4]), .CK(REF_CLK_c), .Q(n7344));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3032 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3030  (.D(n7322[3]), .CK(REF_CLK_c), .Q(n7342));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3030 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3028  (.D(n7322[2]), .CK(REF_CLK_c), .Q(n7340));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3028 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3026  (.D(n7322[1]), .CK(REF_CLK_c), .Q(n7338));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3026 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2972  (.D(n7190[8]), .CK(REF_CLK_c), .Q(n7220));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2972 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3024  (.D(n7322[0]), .CK(REF_CLK_c), .Q(n7336));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3024 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_adj_420  (.D(dmem_write_data[15]), .CK(REF_CLK_c), 
            .Q(n7309));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_adj_420 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3020  (.D(dmem_write_data[14]), .CK(REF_CLK_c), 
            .Q(n7307));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3020 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3019  (.D(dmem_write_data[13]), .CK(REF_CLK_c), 
            .Q(n7305));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3019 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3018  (.D(dmem_write_data[12]), .CK(REF_CLK_c), 
            .Q(n7303));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3018 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3017  (.D(dmem_write_data[11]), .CK(REF_CLK_c), 
            .Q(n7301));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3017 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2970  (.D(n7190[7]), .CK(REF_CLK_c), .Q(n7218));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2970 .GSR = "ENABLED";
    LUT4 mux_3054_i7_3_lut_4_lut (.A(n7358), .B(n7357), .C(n7373), .D(n7372), 
         .Z(n6417[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3054_i7_3_lut_4_lut.init = 16'hf780;
    FD1S3AX \genblk1.mem_3016  (.D(dmem_write_data[10]), .CK(REF_CLK_c), 
            .Q(n7299));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3016 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3015  (.D(dmem_write_data[9]), .CK(REF_CLK_c), 
            .Q(n7297));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3015 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3014  (.D(dmem_write_data[8]), .CK(REF_CLK_c), 
            .Q(n7295));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3014 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3013  (.D(\genblk1.mem_N_2584_adj_179 ), .CK(REF_CLK_c), 
            .Q(n7292));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3013 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3011  (.D(n7256[10]), .CK(REF_CLK_c), .Q(n7290));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3011 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3008  (.D(n7256[9]), .CK(REF_CLK_c), .Q(n7288));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3008 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3006  (.D(n7256[8]), .CK(REF_CLK_c), .Q(n7286));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3006 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3004  (.D(n7256[7]), .CK(REF_CLK_c), .Q(n7284));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3004 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2968  (.D(n7190[6]), .CK(REF_CLK_c), .Q(n7216));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2968 .GSR = "ENABLED";
    LUT4 mux_3054_i8_3_lut_4_lut (.A(n7358), .B(n7357), .C(n7375), .D(n7374), 
         .Z(n6417[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3054_i8_3_lut_4_lut.init = 16'hf780;
    FD1S3AX \genblk1.mem_3002  (.D(n7256[6]), .CK(REF_CLK_c), .Q(n7282));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3002 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_adj_421  (.D(dmem_write_data[31]), .CK(REF_CLK_c), 
            .Q(n7441));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_adj_421 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3088  (.D(dmem_write_data[30]), .CK(REF_CLK_c), 
            .Q(n7439));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3088 .GSR = "ENABLED";
    LUT4 mux_3020_i1_3_lut_4_lut (.A(n7292), .B(n7291), .C(n7295), .D(n7294), 
         .Z(n6416[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3020_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3020_i2_3_lut_4_lut (.A(n7292), .B(n7291), .C(n7297), .D(n7296), 
         .Z(n6416[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3020_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3020_i3_3_lut_4_lut (.A(n7292), .B(n7291), .C(n7299), .D(n7298), 
         .Z(n6416[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3020_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3020_i4_3_lut_4_lut (.A(n7292), .B(n7291), .C(n7301), .D(n7300), 
         .Z(n6416[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3020_i4_3_lut_4_lut.init = 16'hf780;
    FD1S3AX \genblk1.mem_3087  (.D(dmem_write_data[29]), .CK(REF_CLK_c), 
            .Q(n7437));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3087 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3000  (.D(n7256[5]), .CK(REF_CLK_c), .Q(n7280));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3000 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2998  (.D(n7256[4]), .CK(REF_CLK_c), .Q(n7278));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2998 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3086  (.D(dmem_write_data[28]), .CK(REF_CLK_c), 
            .Q(n7435));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3086 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3085  (.D(dmem_write_data[27]), .CK(REF_CLK_c), 
            .Q(n7433));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3085 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2966  (.D(n7190[5]), .CK(REF_CLK_c), .Q(n7214));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2966 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3084  (.D(dmem_write_data[26]), .CK(REF_CLK_c), 
            .Q(n7431));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3084 .GSR = "ENABLED";
    LUT4 mux_3020_i5_3_lut_4_lut (.A(n7292), .B(n7291), .C(n7303), .D(n7302), 
         .Z(n6416[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3020_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3020_i6_3_lut_4_lut (.A(n7292), .B(n7291), .C(n7305), .D(n7304), 
         .Z(n6416[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3020_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3020_i7_3_lut_4_lut (.A(n7292), .B(n7291), .C(n7307), .D(n7306), 
         .Z(n6416[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3020_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3020_i8_3_lut_4_lut (.A(n7292), .B(n7291), .C(n7309), .D(n7308), 
         .Z(n6416[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3020_i8_3_lut_4_lut.init = 16'hf780;
    FD1S3AX \genblk1.mem_2996  (.D(n7256[3]), .CK(REF_CLK_c), .Q(n7276));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2996 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2994  (.D(n7256[2]), .CK(REF_CLK_c), .Q(n7274));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2994 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2992  (.D(n7256[1]), .CK(REF_CLK_c), .Q(n7272));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2992 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3083  (.D(dmem_write_data[25]), .CK(REF_CLK_c), 
            .Q(n7429));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3083 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2965  (.D(dmem_write_address[5]), .CK(REF_CLK_c), 
            .Q(n7279));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_2965 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3082  (.D(dmem_write_data[24]), .CK(REF_CLK_c), 
            .Q(n7427));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3082 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3081  (.D(\genblk1.mem_N_2584_adj_180 ), .CK(REF_CLK_c), 
            .Q(n7424));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3081 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2964  (.D(n7190[4]), .CK(REF_CLK_c), .Q(n7212));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2964 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2963  (.D(dmem_write_address[4]), .CK(REF_CLK_c), 
            .Q(n7277));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_2963 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2990  (.D(n7256[0]), .CK(REF_CLK_c), .Q(n7270));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2990 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3079  (.D(n7388[10]), .CK(REF_CLK_c), .Q(\genblk1.ra [10]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3079 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3076  (.D(n7388[9]), .CK(REF_CLK_c), .Q(\genblk1.ra [9]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3076 .GSR = "ENABLED";
    DP16KD \genblk1.mem0  (.DIA0(dmem_write_data[0]), .DIA1(dmem_write_data[1]), 
           .DIA2(dmem_write_data[2]), .DIA3(dmem_write_data[3]), .DIA4(dmem_write_data[4]), 
           .DIA5(dmem_write_data[5]), .DIA6(dmem_write_data[6]), .DIA7(dmem_write_data[7]), 
           .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), .DIA11(GND_net), 
           .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), .DIA15(GND_net), 
           .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), .ADA1(GND_net), 
           .ADA2(GND_net), .ADA3(dmem_write_address[0]), .ADA4(dmem_write_address[1]), 
           .ADA5(dmem_write_address[2]), .ADA6(dmem_write_address[3]), .ADA7(dmem_write_address[4]), 
           .ADA8(dmem_write_address[5]), .ADA9(dmem_write_address[6]), .ADA10(dmem_write_address[7]), 
           .ADA11(dmem_write_address[8]), .ADA12(dmem_write_address[9]), 
           .ADA13(dmem_write_address[10]), .CEA(VCC_net), .OCEA(VCC_net), 
           .CLKA(REF_CLK_c), .WEA(\genblk1.mem_N_2584_c ), .CSA0(GND_net), 
           .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), 
           .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
           .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
           .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), .DIB12(GND_net), 
           .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), .DIB16(GND_net), 
           .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), 
           .ADB3(n7190[0]), .ADB4(n7190[1]), .ADB5(n7190[2]), .ADB6(n7190[3]), 
           .ADB7(n7190[4]), .ADB8(n7190[5]), .ADB9(n7190[6]), .ADB10(n7190[7]), 
           .ADB11(n7190[8]), .ADB12(n7190[9]), .ADB13(n7190[10]), .CEB(VCC_net), 
           .OCEB(VCC_net), .CLKB(REF_CLK_c), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(GND_net), .DOB0(n7228), 
           .DOB1(n7230), .DOB2(n7232), .DOB3(n7234), .DOB4(n7236), .DOB5(n7238), 
           .DOB6(n7240), .DOB7(n7242));
    defparam \genblk1.mem0 .DATA_WIDTH_A = 9;
    defparam \genblk1.mem0 .DATA_WIDTH_B = 9;
    defparam \genblk1.mem0 .REGMODE_A = "NOREG";
    defparam \genblk1.mem0 .REGMODE_B = "NOREG";
    defparam \genblk1.mem0 .RESETMODE = "SYNC";
    defparam \genblk1.mem0 .ASYNC_RESET_RELEASE = "SYNC";
    defparam \genblk1.mem0 .WRITEMODE_A = "WRITETHROUGH";
    defparam \genblk1.mem0 .WRITEMODE_B = "WRITETHROUGH";
    defparam \genblk1.mem0 .CSDECODE_A = "0b000";
    defparam \genblk1.mem0 .CSDECODE_B = "0b000";
    defparam \genblk1.mem0 .GSR = "DISABLED";
    defparam \genblk1.mem0 .INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INIT_DATA = "STATIC";
    FD1S3AX \genblk1.mem_adj_422  (.D(dmem_write_data[7]), .CK(REF_CLK_c), 
            .Q(n7243));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_adj_422 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3074  (.D(n7388[8]), .CK(REF_CLK_c), .Q(\genblk1.ra [8]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3074 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2962  (.D(n7190[3]), .CK(REF_CLK_c), .Q(n7210));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2962 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3072  (.D(n7388[7]), .CK(REF_CLK_c), .Q(\genblk1.ra [7]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3072 .GSR = "ENABLED";
    CCU2C equal_3077_11 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27381), 
          .S0(n7423));
    defparam equal_3077_11.INIT0 = 16'h0000;
    defparam equal_3077_11.INIT1 = 16'h0000;
    defparam equal_3077_11.INJECT1_0 = "NO";
    defparam equal_3077_11.INJECT1_1 = "NO";
    FD1S3AX \genblk1.mem_2961  (.D(dmem_write_address[3]), .CK(REF_CLK_c), 
            .Q(n7275));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_2961 .GSR = "ENABLED";
    CCU2C equal_3077_11_22479 (.A0(\genblk1.ra [3]), .B0(n7275), .C0(\genblk1.ra [2]), 
          .D0(n7339), .A1(\genblk1.ra [1]), .B1(n7337), .C1(\genblk1.ra [0]), 
          .D1(n7335), .CIN(n27380), .COUT(n27381));
    defparam equal_3077_11_22479.INIT0 = 16'h9009;
    defparam equal_3077_11_22479.INIT1 = 16'h9009;
    defparam equal_3077_11_22479.INJECT1_0 = "YES";
    defparam equal_3077_11_22479.INJECT1_1 = "YES";
    LUT4 i2_4_lut (.A(\byte_enable_m[0] ), .B(n9291), .C(\state[2] ), 
         .D(dcache_select_m), .Z(\genblk1.mem_N_2584_c )) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(298[13:63])
    defparam i2_4_lut.init = 16'hc8c0;
    CCU2C equal_3077_9 (.A0(\genblk1.ra [7]), .B0(n7217), .C0(\genblk1.ra [6]), 
          .D0(n7215), .A1(\genblk1.ra [5]), .B1(n7279), .C1(\genblk1.ra [4]), 
          .D1(n7277), .CIN(n27379), .COUT(n27380));
    defparam equal_3077_9.INIT0 = 16'h9009;
    defparam equal_3077_9.INIT1 = 16'h9009;
    defparam equal_3077_9.INJECT1_0 = "YES";
    defparam equal_3077_9.INJECT1_1 = "YES";
    CCU2C equal_3077_0 (.A0(\genblk1.ra [10]), .B0(n7289), .C0(GND_net), 
          .D0(VCC_net), .A1(\genblk1.ra [9]), .B1(n7287), .C1(\genblk1.ra [8]), 
          .D1(n7285), .COUT(n27379));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam equal_3077_0.INIT0 = 16'h0009;
    defparam equal_3077_0.INIT1 = 16'h9009;
    defparam equal_3077_0.INJECT1_0 = "NO";
    defparam equal_3077_0.INJECT1_1 = "YES";
    CCU2C equal_3009_11 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27378), 
          .S0(n7291));
    defparam equal_3009_11.INIT0 = 16'h0000;
    defparam equal_3009_11.INIT1 = 16'h0000;
    defparam equal_3009_11.INJECT1_0 = "NO";
    defparam equal_3009_11.INJECT1_1 = "NO";
    CCU2C equal_3009_11_22478 (.A0(n7276), .B0(n7275), .C0(n7274), .D0(n7339), 
          .A1(n7272), .B1(n7337), .C1(n7270), .D1(n7335), .CIN(n27377), 
          .COUT(n27378));
    defparam equal_3009_11_22478.INIT0 = 16'h9009;
    defparam equal_3009_11_22478.INIT1 = 16'h9009;
    defparam equal_3009_11_22478.INJECT1_0 = "YES";
    defparam equal_3009_11_22478.INJECT1_1 = "YES";
    CCU2C equal_3009_9 (.A0(n7284), .B0(n7217), .C0(n7282), .D0(n7215), 
          .A1(n7280), .B1(n7279), .C1(n7278), .D1(n7277), .CIN(n27376), 
          .COUT(n27377));
    defparam equal_3009_9.INIT0 = 16'h9009;
    defparam equal_3009_9.INIT1 = 16'h9009;
    defparam equal_3009_9.INJECT1_0 = "YES";
    defparam equal_3009_9.INJECT1_1 = "YES";
    CCU2C equal_3009_0 (.A0(n7290), .B0(n7289), .C0(GND_net), .D0(VCC_net), 
          .A1(n7288), .B1(n7287), .C1(n7286), .D1(n7285), .COUT(n27376));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam equal_3009_0.INIT0 = 16'h0009;
    defparam equal_3009_0.INIT1 = 16'h9009;
    defparam equal_3009_0.INJECT1_0 = "NO";
    defparam equal_3009_0.INJECT1_1 = "YES";
    LUT4 mux_2986_i1_3_lut_4_lut (.A(n7226), .B(n7225), .C(n7229), .D(n7228), 
         .Z(dcache_data_m[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_2986_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_2986_i2_3_lut_4_lut (.A(n7226), .B(n7225), .C(n7231), .D(n7230), 
         .Z(dcache_data_m[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_2986_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_2986_i3_3_lut_4_lut (.A(n7226), .B(n7225), .C(n7233), .D(n7232), 
         .Z(dcache_data_m[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_2986_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_2986_i4_3_lut_4_lut (.A(n7226), .B(n7225), .C(n7235), .D(n7234), 
         .Z(dcache_data_m[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_2986_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_2986_i5_3_lut_4_lut (.A(n7226), .B(n7225), .C(n7237), .D(n7236), 
         .Z(dcache_data_m[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_2986_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_2986_i6_3_lut_4_lut (.A(n7226), .B(n7225), .C(n7239), .D(n7238), 
         .Z(dcache_data_m[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_2986_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_2986_i7_3_lut_4_lut (.A(n7226), .B(n7225), .C(n7241), .D(n7240), 
         .Z(dcache_data_m[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_2986_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_2986_i8_3_lut_4_lut (.A(n7226), .B(n7225), .C(n7243), .D(n7242), 
         .Z(dcache_data_m[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_2986_i8_3_lut_4_lut.init = 16'hf780;
    CCU2C equal_3043_11 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27371), 
          .S0(n7357));
    defparam equal_3043_11.INIT0 = 16'h0000;
    defparam equal_3043_11.INIT1 = 16'h0000;
    defparam equal_3043_11.INJECT1_0 = "NO";
    defparam equal_3043_11.INJECT1_1 = "NO";
    CCU2C equal_3043_11_22477 (.A0(n7342), .B0(n7275), .C0(n7340), .D0(n7339), 
          .A1(n7338), .B1(n7337), .C1(n7336), .D1(n7335), .CIN(n27370), 
          .COUT(n27371));
    defparam equal_3043_11_22477.INIT0 = 16'h9009;
    defparam equal_3043_11_22477.INIT1 = 16'h9009;
    defparam equal_3043_11_22477.INJECT1_0 = "YES";
    defparam equal_3043_11_22477.INJECT1_1 = "YES";
    CCU2C equal_3043_9 (.A0(n7350), .B0(n7217), .C0(n7348), .D0(n7215), 
          .A1(n7346), .B1(n7279), .C1(n7344), .D1(n7277), .CIN(n27369), 
          .COUT(n27370));
    defparam equal_3043_9.INIT0 = 16'h9009;
    defparam equal_3043_9.INIT1 = 16'h9009;
    defparam equal_3043_9.INJECT1_0 = "YES";
    defparam equal_3043_9.INJECT1_1 = "YES";
    CCU2C equal_3043_0 (.A0(n7356), .B0(n7289), .C0(GND_net), .D0(VCC_net), 
          .A1(n7354), .B1(n7287), .C1(n7352), .D1(n7285), .COUT(n27369));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam equal_3043_0.INIT0 = 16'h0009;
    defparam equal_3043_0.INIT1 = 16'h9009;
    defparam equal_3043_0.INJECT1_0 = "NO";
    defparam equal_3043_0.INJECT1_1 = "YES";
    CCU2C equal_2975_11 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27368), 
          .S0(n7225));
    defparam equal_2975_11.INIT0 = 16'h0000;
    defparam equal_2975_11.INIT1 = 16'h0000;
    defparam equal_2975_11.INJECT1_0 = "NO";
    defparam equal_2975_11.INJECT1_1 = "NO";
    CCU2C equal_2975_11_22476 (.A0(n7210), .B0(n7275), .C0(n7208), .D0(n7339), 
          .A1(n7206), .B1(n7337), .C1(n7204), .D1(n7335), .CIN(n27367), 
          .COUT(n27368));
    defparam equal_2975_11_22476.INIT0 = 16'h9009;
    defparam equal_2975_11_22476.INIT1 = 16'h9009;
    defparam equal_2975_11_22476.INJECT1_0 = "YES";
    defparam equal_2975_11_22476.INJECT1_1 = "YES";
    CCU2C equal_2975_9 (.A0(n7218), .B0(n7217), .C0(n7216), .D0(n7215), 
          .A1(n7214), .B1(n7279), .C1(n7212), .D1(n7277), .CIN(n27366), 
          .COUT(n27367));
    defparam equal_2975_9.INIT0 = 16'h9009;
    defparam equal_2975_9.INIT1 = 16'h9009;
    defparam equal_2975_9.INJECT1_0 = "YES";
    defparam equal_2975_9.INJECT1_1 = "YES";
    
endmodule
//
// Verilog Description of module lm32_jtag
//

module lm32_jtag (jtag_reg_q, jtag_reg_d_7__N_515, jtag_reg_d, REF_CLK_c, 
            REF_CLK_c_enable_1373, REF_CLK_c_enable_1606, n4626, rx_toggle_r_r, 
            rx_toggle_r_r_r, uart_tx_byte, \operand_1_x[0] , \jrx_csr_read_data[0] , 
            jrx_csr_read_data_8__N_3304, jtag_break, reset_exception, 
            \jtag_reg_addr_d[0] , \jtag_reg_addr_d[1] , jtag_update_N_3371, 
            \operand_1_x[1] , \operand_1_x[2] , \operand_1_x[3] , \operand_1_x[4] , 
            \operand_1_x[5] , \operand_1_x[6] , \operand_1_x[7] , \jrx_csr_read_data[1] , 
            \jrx_csr_read_data[2] , \jrx_csr_read_data[3] , \jrx_csr_read_data[4] , 
            \jrx_csr_read_data[5] , \jrx_csr_read_data[6] , \jrx_csr_read_data[7] , 
            n41232, n4, n41233, n34542, \jtag_reg_addr_q[1] , n30162, 
            n43, n33932, n29834, n34464) /* synthesis syn_module_defined=1 */ ;
    input [7:0]jtag_reg_q;
    input jtag_reg_d_7__N_515;
    output [7:0]jtag_reg_d;
    input REF_CLK_c;
    input REF_CLK_c_enable_1373;
    input REF_CLK_c_enable_1606;
    input [7:0]n4626;
    output rx_toggle_r_r;
    output rx_toggle_r_r_r;
    output [7:0]uart_tx_byte;
    input \operand_1_x[0] ;
    output \jrx_csr_read_data[0] ;
    input jrx_csr_read_data_8__N_3304;
    output jtag_break;
    output reset_exception;
    output \jtag_reg_addr_d[0] ;
    output \jtag_reg_addr_d[1] ;
    input jtag_update_N_3371;
    input \operand_1_x[1] ;
    input \operand_1_x[2] ;
    input \operand_1_x[3] ;
    input \operand_1_x[4] ;
    input \operand_1_x[5] ;
    input \operand_1_x[6] ;
    input \operand_1_x[7] ;
    output \jrx_csr_read_data[1] ;
    output \jrx_csr_read_data[2] ;
    output \jrx_csr_read_data[3] ;
    output \jrx_csr_read_data[4] ;
    output \jrx_csr_read_data[5] ;
    output \jrx_csr_read_data[6] ;
    output \jrx_csr_read_data[7] ;
    input n41232;
    input n4;
    input n41233;
    input n34542;
    input \jtag_reg_addr_q[1] ;
    input n30162;
    input n43;
    input n33932;
    input n29834;
    input n34464;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire jtag_update_N_3371 /* synthesis is_inv_clock=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(203[14:23])
    
    wire n29798, n41211, REF_CLK_c_enable_169, n41212, REF_CLK_c_enable_168, 
        rx_toggle_r, rx_toggle, REF_CLK_c_enable_1409, jtx_csr_read_data_8__N_3287, 
        REF_CLK_c_enable_170, rx_toggle_N_3369, n30163;
    
    LUT4 i33142_2_lut_rep_806 (.A(jtag_reg_q[4]), .B(n29798), .Z(n41211)) /* synthesis lut_function=(!((B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(429[7:15])
    defparam i33142_2_lut_rep_806.init = 16'h2222;
    LUT4 i1_2_lut_3_lut (.A(jtag_reg_q[4]), .B(n29798), .C(jtag_reg_d_7__N_515), 
         .Z(REF_CLK_c_enable_169)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(429[7:15])
    defparam i1_2_lut_3_lut.init = 16'hf2f2;
    LUT4 i33145_2_lut_rep_807 (.A(jtag_reg_q[4]), .B(n29798), .Z(n41212)) /* synthesis lut_function=(!(A+(B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(450[7:21])
    defparam i33145_2_lut_rep_807.init = 16'h1111;
    LUT4 i1_2_lut_3_lut_adj_417 (.A(jtag_reg_q[4]), .B(n29798), .C(jtag_reg_d_7__N_515), 
         .Z(REF_CLK_c_enable_168)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(450[7:21])
    defparam i1_2_lut_3_lut_adj_417.init = 16'hf1f1;
    FD1P3DX jtag_reg_d_i0_i0 (.D(n4626[0]), .SP(REF_CLK_c_enable_1373), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(jtag_reg_d[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reg_d_i0_i0.GSR = "ENABLED";
    FD1S3DX rx_toggle_r_82 (.D(rx_toggle), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(rx_toggle_r)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(301[4] 305[7])
    defparam rx_toggle_r_82.GSR = "ENABLED";
    FD1S3DX rx_toggle_r_r_83 (.D(rx_toggle_r), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(rx_toggle_r_r)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(301[4] 305[7])
    defparam rx_toggle_r_r_83.GSR = "ENABLED";
    FD1S3DX rx_toggle_r_r_r_84 (.D(rx_toggle_r_r), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(rx_toggle_r_r_r)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(301[4] 305[7])
    defparam rx_toggle_r_r_r_84.GSR = "ENABLED";
    FD1P3DX uart_tx_byte_i0_i0 (.D(\operand_1_x[0] ), .SP(REF_CLK_c_enable_1409), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(uart_tx_byte[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_byte_i0_i0.GSR = "ENABLED";
    FD1P3DX uart_rx_byte__i1 (.D(jtag_reg_q[0]), .SP(jrx_csr_read_data_8__N_3304), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\jrx_csr_read_data[0] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_byte__i1.GSR = "ENABLED";
    FD1P3DX jtag_break_88 (.D(n41212), .SP(REF_CLK_c_enable_168), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(jtag_break)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_break_88.GSR = "ENABLED";
    FD1P3DX jtag_reset_89 (.D(n41211), .SP(REF_CLK_c_enable_169), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reset_exception)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reset_89.GSR = "ENABLED";
    FD1S3DX uart_tx_valid_91 (.D(jtx_csr_read_data_8__N_3287), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\jtag_reg_addr_d[0] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_valid_91.GSR = "ENABLED";
    FD1P3DX uart_rx_valid_93 (.D(jrx_csr_read_data_8__N_3304), .SP(REF_CLK_c_enable_170), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\jtag_reg_addr_d[1] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_valid_93.GSR = "ENABLED";
    FD1S3DX rx_toggle_81 (.D(rx_toggle_N_3369), .CK(jtag_update_N_3371), 
            .CD(REF_CLK_c_enable_1606), .Q(rx_toggle)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(279[4:31])
    defparam rx_toggle_81.GSR = "ENABLED";
    FD1P3DX jtag_reg_d_i0_i1 (.D(n4626[1]), .SP(REF_CLK_c_enable_1373), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(jtag_reg_d[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reg_d_i0_i1.GSR = "ENABLED";
    FD1P3DX jtag_reg_d_i0_i2 (.D(n4626[2]), .SP(REF_CLK_c_enable_1373), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(jtag_reg_d[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reg_d_i0_i2.GSR = "ENABLED";
    FD1P3DX jtag_reg_d_i0_i3 (.D(n4626[3]), .SP(REF_CLK_c_enable_1373), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(jtag_reg_d[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reg_d_i0_i3.GSR = "ENABLED";
    FD1P3DX jtag_reg_d_i0_i4 (.D(n4626[4]), .SP(REF_CLK_c_enable_1373), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(jtag_reg_d[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reg_d_i0_i4.GSR = "ENABLED";
    FD1P3DX jtag_reg_d_i0_i5 (.D(n4626[5]), .SP(REF_CLK_c_enable_1373), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(jtag_reg_d[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reg_d_i0_i5.GSR = "ENABLED";
    FD1P3DX jtag_reg_d_i0_i6 (.D(n4626[6]), .SP(REF_CLK_c_enable_1373), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(jtag_reg_d[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reg_d_i0_i6.GSR = "ENABLED";
    FD1P3DX jtag_reg_d_i0_i7 (.D(n4626[7]), .SP(REF_CLK_c_enable_1373), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(jtag_reg_d[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reg_d_i0_i7.GSR = "ENABLED";
    FD1P3DX uart_tx_byte_i0_i1 (.D(\operand_1_x[1] ), .SP(REF_CLK_c_enable_1409), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(uart_tx_byte[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_byte_i0_i1.GSR = "ENABLED";
    FD1P3DX uart_tx_byte_i0_i2 (.D(\operand_1_x[2] ), .SP(REF_CLK_c_enable_1409), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(uart_tx_byte[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_byte_i0_i2.GSR = "ENABLED";
    FD1P3DX uart_tx_byte_i0_i3 (.D(\operand_1_x[3] ), .SP(REF_CLK_c_enable_1409), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(uart_tx_byte[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_byte_i0_i3.GSR = "ENABLED";
    FD1P3DX uart_tx_byte_i0_i4 (.D(\operand_1_x[4] ), .SP(REF_CLK_c_enable_1409), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(uart_tx_byte[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_byte_i0_i4.GSR = "ENABLED";
    FD1P3DX uart_tx_byte_i0_i5 (.D(\operand_1_x[5] ), .SP(REF_CLK_c_enable_1409), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(uart_tx_byte[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_byte_i0_i5.GSR = "ENABLED";
    FD1P3DX uart_tx_byte_i0_i6 (.D(\operand_1_x[6] ), .SP(REF_CLK_c_enable_1409), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(uart_tx_byte[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_byte_i0_i6.GSR = "ENABLED";
    FD1P3DX uart_tx_byte_i0_i7 (.D(\operand_1_x[7] ), .SP(REF_CLK_c_enable_1409), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(uart_tx_byte[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_byte_i0_i7.GSR = "ENABLED";
    FD1P3DX uart_rx_byte__i2 (.D(jtag_reg_q[1]), .SP(jrx_csr_read_data_8__N_3304), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\jrx_csr_read_data[1] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_byte__i2.GSR = "ENABLED";
    FD1P3DX uart_rx_byte__i3 (.D(jtag_reg_q[2]), .SP(jrx_csr_read_data_8__N_3304), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\jrx_csr_read_data[2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_byte__i3.GSR = "ENABLED";
    FD1P3DX uart_rx_byte__i4 (.D(jtag_reg_q[3]), .SP(jrx_csr_read_data_8__N_3304), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\jrx_csr_read_data[3] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_byte__i4.GSR = "ENABLED";
    FD1P3DX uart_rx_byte__i5 (.D(jtag_reg_q[4]), .SP(jrx_csr_read_data_8__N_3304), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\jrx_csr_read_data[4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_byte__i5.GSR = "ENABLED";
    FD1P3DX uart_rx_byte__i6 (.D(jtag_reg_q[5]), .SP(jrx_csr_read_data_8__N_3304), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\jrx_csr_read_data[5] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_byte__i6.GSR = "ENABLED";
    FD1P3DX uart_rx_byte__i7 (.D(jtag_reg_q[6]), .SP(jrx_csr_read_data_8__N_3304), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\jrx_csr_read_data[6] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_byte__i7.GSR = "ENABLED";
    FD1P3DX uart_rx_byte__i8 (.D(jtag_reg_q[7]), .SP(jrx_csr_read_data_8__N_3304), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\jrx_csr_read_data[7] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_byte__i8.GSR = "ENABLED";
    LUT4 i33147_4_lut (.A(n41232), .B(n4), .C(n41233), .D(n34542), .Z(REF_CLK_c_enable_1409)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i33147_4_lut.init = 16'h0008;
    LUT4 i1_4_lut (.A(\jtag_reg_addr_q[1] ), .B(n30162), .C(jtag_reg_q[7]), 
         .D(n43), .Z(n29798)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(427[5] 493[12])
    defparam i1_4_lut.init = 16'hfeff;
    LUT4 i14639_4_lut (.A(\jtag_reg_addr_d[0] ), .B(n30163), .C(n33932), 
         .D(n4), .Z(jtx_csr_read_data_8__N_3287)) /* synthesis lut_function=(A (B)+!A !((C+!(D))+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(424[7] 494[12])
    defparam i14639_4_lut.init = 16'h8c88;
    LUT4 i1_4_lut_adj_418 (.A(jtag_reg_q[7]), .B(n30162), .C(\jtag_reg_addr_q[1] ), 
         .D(n43), .Z(n30163)) /* synthesis lut_function=(A (B+!(C))+!A (B+!(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(424[7] 494[12])
    defparam i1_4_lut_adj_418.init = 16'hcecf;
    LUT4 i1_4_lut_adj_419 (.A(n41232), .B(n29834), .C(n4), .D(n34464), 
         .Z(REF_CLK_c_enable_170)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut_adj_419.init = 16'hccec;
    LUT4 rx_toggle_I_0_1_lut (.A(rx_toggle), .Z(rx_toggle_N_3369)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(279[20:30])
    defparam rx_toggle_I_0_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module lm32_interrupt
//

module lm32_interrupt (csr_x, n41288, im, REF_CLK_c, REF_CLK_c_enable_1335, 
            REF_CLK_c_enable_1606, operand_1_x, n41308, n4354, bie, 
            REF_CLK_c_enable_391, n36337, n9401, ie, \im[2] , \im[3] , 
            \im[4] , \im[5] , \im[6] , \im[7] , \im[8] , \im[9] , 
            \im[10] , \im[11] , \im[12] , \im[13] , \im[14] , \im[15] , 
            \im[16] , \im[17] , \im[18] , \im[19] , \im[20] , \im[21] , 
            \im[22] , \im[23] , \im[24] , \im[25] , \im[26] , \im[27] , 
            \im[28] , \im[29] , \im[30] , \im[31] , \ip[1] , n32134, 
            store_x, n32132, n41313, n41393, n41391, n31825, n11934, 
            n45175, branch_flushX_m, n35639, dcache_refill_request, 
            n35022, eret_q_x, n34986, n35030, valid_w, non_debug_exception_w, 
            debug_exception_w, n41240, n41394, eret_x, bret_x, n41400, 
            n34542, valid_x, n20581, n41232, n34942, SPI_INT_O_N_4422, 
            SPI_INT_O_N_4417, SPI_INT_O_N_4421, n31334, n41183, n41401, 
            n41317, n41413, n34898, n41416, LM32D_CYC_O, n33946) /* synthesis syn_module_defined=1 */ ;
    input [4:0]csr_x;
    output n41288;
    output [31:0]im;
    input REF_CLK_c;
    input REF_CLK_c_enable_1335;
    input REF_CLK_c_enable_1606;
    input [31:0]operand_1_x;
    output n41308;
    output n4354;
    output bie;
    input REF_CLK_c_enable_391;
    input n36337;
    input n9401;
    output ie;
    output \im[2] ;
    output \im[3] ;
    output \im[4] ;
    output \im[5] ;
    output \im[6] ;
    output \im[7] ;
    output \im[8] ;
    output \im[9] ;
    output \im[10] ;
    output \im[11] ;
    output \im[12] ;
    output \im[13] ;
    output \im[14] ;
    output \im[15] ;
    output \im[16] ;
    output \im[17] ;
    output \im[18] ;
    output \im[19] ;
    output \im[20] ;
    output \im[21] ;
    output \im[22] ;
    output \im[23] ;
    output \im[24] ;
    output \im[25] ;
    output \im[26] ;
    output \im[27] ;
    output \im[28] ;
    output \im[29] ;
    output \im[30] ;
    output \im[31] ;
    output \ip[1] ;
    output n32134;
    input store_x;
    output n32132;
    output n41313;
    output n41393;
    input n41391;
    output n31825;
    output n11934;
    input n45175;
    input branch_flushX_m;
    output n35639;
    input dcache_refill_request;
    input n35022;
    input eret_q_x;
    input n34986;
    input n35030;
    input valid_w;
    input non_debug_exception_w;
    input debug_exception_w;
    output n41240;
    output n41394;
    input eret_x;
    input bret_x;
    output n41400;
    output n34542;
    input valid_x;
    input n20581;
    input n41232;
    input n34942;
    input SPI_INT_O_N_4422;
    input SPI_INT_O_N_4417;
    input SPI_INT_O_N_4421;
    input n31334;
    input n41183;
    input n41401;
    output n41317;
    input n41413;
    output n34898;
    output n41416;
    input LM32D_CYC_O;
    output n33946;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    
    wire n41412, eie;
    wire [31:0]im_c;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(141[22:24])
    
    wire REF_CLK_c_enable_392, REF_CLK_c_enable_1233, n12407;
    wire [31:0]ip_31__N_3128;
    
    wire n35765, n41314, ie_N_3261;
    wire [31:0]asserted;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(129[23:31])
    
    wire n35932, n35786;
    
    LUT4 i1_2_lut_rep_883_4_lut (.A(csr_x[2]), .B(n41412), .C(csr_x[1]), 
         .D(csr_x[0]), .Z(n41288)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_883_4_lut.init = 16'h0100;
    FD1P3DX im_i0_i0 (.D(operand_1_x[0]), .SP(REF_CLK_c_enable_1335), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(im[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i0.GSR = "ENABLED";
    LUT4 i14927_4_lut (.A(eie), .B(n41308), .C(im_c[1]), .D(csr_x[0]), 
         .Z(n4354)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(173[5] 186[12])
    defparam i14927_4_lut.init = 16'h3022;
    FD1P3DX bie_68 (.D(n36337), .SP(REF_CLK_c_enable_391), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(bie)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam bie_68.GSR = "ENABLED";
    FD1P3DX eie_67 (.D(n9401), .SP(REF_CLK_c_enable_392), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(eie)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam eie_67.GSR = "ENABLED";
    FD1P3DX ie_66 (.D(n12407), .SP(REF_CLK_c_enable_1233), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(ie)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam ie_66.GSR = "ENABLED";
    FD1P3DX im_i0_i1 (.D(operand_1_x[1]), .SP(REF_CLK_c_enable_1335), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(im_c[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i1.GSR = "ENABLED";
    FD1P3DX im_i0_i2 (.D(operand_1_x[2]), .SP(REF_CLK_c_enable_1335), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\im[2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i2.GSR = "ENABLED";
    FD1P3DX im_i0_i3 (.D(operand_1_x[3]), .SP(REF_CLK_c_enable_1335), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\im[3] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i3.GSR = "ENABLED";
    FD1P3DX im_i0_i4 (.D(operand_1_x[4]), .SP(REF_CLK_c_enable_1335), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\im[4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i4.GSR = "ENABLED";
    FD1P3DX im_i0_i5 (.D(operand_1_x[5]), .SP(REF_CLK_c_enable_1335), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\im[5] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i5.GSR = "ENABLED";
    FD1P3DX im_i0_i6 (.D(operand_1_x[6]), .SP(REF_CLK_c_enable_1335), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\im[6] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i6.GSR = "ENABLED";
    FD1P3DX im_i0_i7 (.D(operand_1_x[7]), .SP(REF_CLK_c_enable_1335), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\im[7] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i7.GSR = "ENABLED";
    FD1P3DX im_i0_i8 (.D(operand_1_x[8]), .SP(REF_CLK_c_enable_1335), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\im[8] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i8.GSR = "ENABLED";
    FD1P3DX im_i0_i9 (.D(operand_1_x[9]), .SP(REF_CLK_c_enable_1335), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\im[9] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i9.GSR = "ENABLED";
    FD1P3DX im_i0_i10 (.D(operand_1_x[10]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[10] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i10.GSR = "ENABLED";
    FD1P3DX im_i0_i11 (.D(operand_1_x[11]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[11] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i11.GSR = "ENABLED";
    FD1P3DX im_i0_i12 (.D(operand_1_x[12]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[12] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i12.GSR = "ENABLED";
    FD1P3DX im_i0_i13 (.D(operand_1_x[13]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[13] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i13.GSR = "ENABLED";
    FD1P3DX im_i0_i14 (.D(operand_1_x[14]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[14] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i14.GSR = "ENABLED";
    FD1P3DX im_i0_i15 (.D(operand_1_x[15]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[15] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i15.GSR = "ENABLED";
    FD1P3DX im_i0_i16 (.D(operand_1_x[16]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[16] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i16.GSR = "ENABLED";
    FD1P3DX im_i0_i17 (.D(operand_1_x[17]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[17] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i17.GSR = "ENABLED";
    FD1P3DX im_i0_i18 (.D(operand_1_x[18]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[18] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i18.GSR = "ENABLED";
    FD1P3DX im_i0_i19 (.D(operand_1_x[19]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[19] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i19.GSR = "ENABLED";
    FD1P3DX im_i0_i20 (.D(operand_1_x[20]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[20] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i20.GSR = "ENABLED";
    FD1P3DX im_i0_i21 (.D(operand_1_x[21]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[21] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i21.GSR = "ENABLED";
    FD1P3DX im_i0_i22 (.D(operand_1_x[22]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[22] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i22.GSR = "ENABLED";
    FD1P3DX im_i0_i23 (.D(operand_1_x[23]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[23] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i23.GSR = "ENABLED";
    FD1P3DX im_i0_i24 (.D(operand_1_x[24]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[24] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i24.GSR = "ENABLED";
    FD1P3DX im_i0_i25 (.D(operand_1_x[25]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[25] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i25.GSR = "ENABLED";
    FD1P3DX im_i0_i26 (.D(operand_1_x[26]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[26] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i26.GSR = "ENABLED";
    FD1P3DX im_i0_i27 (.D(operand_1_x[27]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[27] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i27.GSR = "ENABLED";
    FD1P3DX im_i0_i28 (.D(operand_1_x[28]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[28] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i28.GSR = "ENABLED";
    FD1P3DX im_i0_i29 (.D(operand_1_x[29]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[29] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i29.GSR = "ENABLED";
    FD1P3DX im_i0_i30 (.D(operand_1_x[30]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[30] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i30.GSR = "ENABLED";
    FD1P3DX im_i0_i31 (.D(operand_1_x[31]), .SP(REF_CLK_c_enable_1335), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\im[31] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i31.GSR = "ENABLED";
    FD1S3DX ip_i1 (.D(ip_31__N_3128[1]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\ip[1] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam ip_i1.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(ie), .B(\ip[1] ), .Z(n32134)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(151[30:59])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_413 (.A(im_c[1]), .B(store_x), .Z(n32132)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(151[30:59])
    defparam i1_2_lut_adj_413.init = 16'h8888;
    LUT4 i33282_3_lut_4_lut (.A(n41313), .B(n41393), .C(n41391), .D(n41308), 
         .Z(n31825)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(183[5:17])
    defparam i33282_3_lut_4_lut.init = 16'h000e;
    LUT4 i7040_4_lut (.A(n11934), .B(n45175), .C(branch_flushX_m), .D(n35765), 
         .Z(REF_CLK_c_enable_1233)) /* synthesis lut_function=(A+!((C+!(D))+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam i7040_4_lut.init = 16'haeaa;
    LUT4 i1_4_lut (.A(n35639), .B(n41314), .C(dcache_refill_request), 
         .D(n35022), .Z(n35765)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;
    defparam i1_4_lut.init = 16'hcdcc;
    LUT4 i14727_4_lut (.A(ie_N_3261), .B(n11934), .C(eie), .D(eret_q_x), 
         .Z(n12407)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam i14727_4_lut.init = 16'h3022;
    LUT4 ie_I_130_4_lut (.A(n34986), .B(bie), .C(n35030), .D(branch_flushX_m), 
         .Z(ie_N_3261)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(266[18] 281[16])
    defparam ie_I_130_4_lut.init = 16'h00ca;
    LUT4 i6582_3_lut (.A(valid_w), .B(non_debug_exception_w), .C(debug_exception_w), 
         .Z(n11934)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i6582_3_lut.init = 16'ha8a8;
    LUT4 i1_2_lut_rep_988 (.A(csr_x[0]), .B(csr_x[1]), .Z(n41393)) /* synthesis lut_function=(A+!(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(183[5:17])
    defparam i1_2_lut_rep_988.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_835_3_lut_4_lut (.A(csr_x[0]), .B(csr_x[1]), .C(csr_x[2]), 
         .D(n41412), .Z(n41240)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(183[5:17])
    defparam i1_2_lut_rep_835_3_lut_4_lut.init = 16'hfffb;
    LUT4 csr_4__I_0_71_i6_2_lut_rep_989 (.A(csr_x[0]), .B(csr_x[1]), .Z(n41394)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(174[5:17])
    defparam csr_4__I_0_71_i6_2_lut_rep_989.init = 16'heeee;
    LUT4 i30481_2_lut_3_lut_4_lut (.A(csr_x[0]), .B(csr_x[1]), .C(csr_x[2]), 
         .D(n41412), .Z(n35639)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(174[5:17])
    defparam i30481_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i15315_2_lut_rep_995 (.A(eret_x), .B(bret_x), .Z(n41400)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i15315_2_lut_rep_995.init = 16'heeee;
    LUT4 i1_4_lut_adj_414 (.A(csr_x[1]), .B(csr_x[3]), .C(csr_x[0]), .D(csr_x[4]), 
         .Z(n34542)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_4_lut_adj_414.init = 16'hfff7;
    LUT4 i1_3_lut_rep_909_4_lut (.A(eret_x), .B(bret_x), .C(valid_x), 
         .D(dcache_refill_request), .Z(n41314)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i1_3_lut_rep_909_4_lut.init = 16'h00e0;
    LUT4 i4567_4_lut (.A(n20581), .B(asserted[1]), .C(n41232), .D(n34942), 
         .Z(ip_31__N_3128[1])) /* synthesis lut_function=(A (B)+!A (B ((D)+!C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(279[17] 280[73])
    defparam i4567_4_lut.init = 16'hcc8c;
    LUT4 i1_4_lut_adj_415 (.A(SPI_INT_O_N_4422), .B(SPI_INT_O_N_4417), .C(SPI_INT_O_N_4421), 
         .D(\ip[1] ), .Z(asserted[1])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(154[19:36])
    defparam i1_4_lut_adj_415.init = 16'hfffe;
    LUT4 i1_4_lut_adj_416 (.A(n31334), .B(REF_CLK_c_enable_391), .C(n41183), 
         .D(n35932), .Z(REF_CLK_c_enable_392)) /* synthesis lut_function=(!(A (B)+!A (B ((D)+!C)))) */ ;
    defparam i1_4_lut_adj_416.init = 16'h3373;
    LUT4 i30770_4_lut (.A(n35786), .B(n41394), .C(n41401), .D(csr_x[3]), 
         .Z(n35932)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30770_4_lut.init = 16'hfffe;
    LUT4 i30624_2_lut (.A(csr_x[2]), .B(csr_x[4]), .Z(n35786)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i30624_2_lut.init = 16'heeee;
    LUT4 equal_1588_i6_2_lut_rep_1007 (.A(csr_x[3]), .B(csr_x[4]), .Z(n41412)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(183[5:17])
    defparam equal_1588_i6_2_lut_rep_1007.init = 16'heeee;
    LUT4 i1_3_lut_rep_903_4_lut (.A(csr_x[3]), .B(csr_x[4]), .C(csr_x[1]), 
         .D(csr_x[2]), .Z(n41308)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(183[5:17])
    defparam i1_3_lut_rep_903_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_912_3_lut (.A(csr_x[3]), .B(csr_x[4]), .C(csr_x[2]), 
         .Z(n41317)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(183[5:17])
    defparam i1_2_lut_rep_912_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_rep_908_3_lut (.A(csr_x[3]), .B(csr_x[4]), .C(csr_x[2]), 
         .Z(n41313)) /* synthesis lut_function=(A+(B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(183[5:17])
    defparam i1_2_lut_rep_908_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(csr_x[3]), .B(csr_x[4]), .C(n41413), 
         .D(csr_x[2]), .Z(n34898)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(183[5:17])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_3_lut_rep_1011 (.A(\ip[1] ), .B(ie), .C(im_c[1]), .Z(n41416)) /* synthesis lut_function=(A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(151[30:59])
    defparam i1_3_lut_rep_1011.init = 16'h8080;
    LUT4 i1_2_lut_4_lut (.A(\ip[1] ), .B(ie), .C(im_c[1]), .D(LM32D_CYC_O), 
         .Z(n33946)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(151[30:59])
    defparam i1_2_lut_4_lut.init = 16'h0080;
    
endmodule
//
// Verilog Description of module \lm32_instruction_unit(base_address=32'b0,limit=32'b01111111111111111) 
//

module \lm32_instruction_unit(base_address=32'b0,limit=32'b01111111111111111)  (\genblk1.wait_one_tick_done , 
            n6781, n41208, n6764, n6769, n6749, REF_CLK_c, stall_a, 
            way_match_0__N_2007, bus_error_f_N_1884, n41410, n13990, 
            n32216, n45075, n41244, n41419, n41295, n41248, n30216, 
            REF_CLK_c_enable_1606, VCC_net, n41178, \LM32I_CTI_O[0] , 
            REF_CLK_c_enable_97, n30900, pc_d, REF_CLK_c_enable_1178, 
            pc_f, pc_x, REF_CLK_c_enable_1624, pc_m, REF_CLK_c_enable_1235, 
            REF_CLK_c_enable_1131, SHAREDBUS_DAT_O, n6760, n6765, n31717, 
            n45105, n6771, n73, n41461, n41228, n41365, n41361, 
            scall_d, n41437, n6778, n6780, n31542, n6768, n32910, 
            n6779, n10, n6777, n6775, branch_taken_m, icache_refill_request, 
            \next_cycle_type[2] , n45080, n41390, n5223, n37955, n37956, 
            n37954, n41345, n41250, n41251, n41279, \LM32I_ADR_O[2] , 
            n45079, \reg_12[2] , n2, \reg_12[12] , n40677, \reg_12[29] , 
            n2_adj_149, \reg_12[3] , n2_adj_150, \reg_12[6] , n2_adj_151, 
            \reg_12[4] , n2_adj_152, \reg_12[14] , n2_adj_153, n30241, 
            n31750, n31955, n41429, \reg_12[22] , n2_adj_154, \reg_12[13] , 
            n2_adj_155, \reg_12[21] , n2_adj_156, \reg_12[28] , n2_adj_157, 
            \reg_12[11] , n2_adj_158, \reg_12[18] , n2_adj_159, \reg_12[25] , 
            n2_adj_160, \reg_12[9] , n2_adj_161, \reg_12[17] , n2_adj_162, 
            \reg_12[24] , n2_adj_163, \reg_12[7] , n2_adj_164, \reg_12[15] , 
            n2_adj_165, n41382, n45183, n6770, n6589, n6584, n37179, 
            \write_idx_x[0] , n35751, n35860, n6439, n6434, n37177, 
            n6599, n6594, n37180, n6629, n6624, n37183, n6579, 
            n6574, n37178, n6429, n6424, n37176, n45103, n35687, 
            n35832, n6609, n6604, n37181, n6619, n6614, n37182, 
            n37185, n37184, n37188, n37187, n37186, n37189, n7603, 
            n7571, n7609, n7607, n7575, n7606, n7574, bus_error_d, 
            n7604, n7572, n7605, n7573, n7608, n7576, n7602, n7570, 
            \selected_1__N_354[0] , n7601, n7569, n7600, n7568, n7599, 
            n7567, n7598, n7566, n7597, n7565, n7596, n7564, n7595, 
            n7563, n7594, n7562, n7593, n7561, n7592, n7560, n7584, 
            n7552, n7583, n7551, n7582, n7550, n7581, n7549, n7580, 
            n7548, n7579, n7547, n7578, n7546, n7577, n7545, n6750, 
            n7591, n7559, n7590, n7558, n7589, n7557, n7588, n7556, 
            n7587, n7555, n7586, n7554, n7585, n7553, n4, \write_idx_x[3] , 
            n32116, n41430, \write_idx_w[3] , n33920, n37501, n37500, 
            n37502, n37499, n37498, n37497, n37496, n6751, n6752, 
            n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6761, 
            n6762, n6763, n6766, n6767, n6776, n40094, n37495, 
            n7672, n7640, n7677, n7673, n7641, \write_idx_x[4] , 
            n32260, n32262, n41312, n41296, n34, n7674, n7642, 
            n7675, n7643, n7676, n7644, n7671, n7639, n7670, n7638, 
            n7669, n7637, n7668, n7636, n7667, n7635, n7666, n7634, 
            n7665, n7633, n7664, n7632, n7663, n7631, n7662, n7630, 
            n7661, n7629, n7660, n7628, n36, n7652, n7620, n7651, 
            n7619, n7650, n7618, n7649, n7617, n37, n7648, n7616, 
            n7647, n7615, n7646, n7614, n7645, n7613, n7659, n7627, 
            n7658, n7626, n7657, n7625, n7656, n7624, n7655, n7623, 
            n7654, n7622, n7653, n7621, n30012, \write_idx_m[2] , 
            n31976, n37504, n37503, n37507, n37506, n37505, n37508, 
            n41364, n41363, n30820, n11834, n41216, n32356, n41281, 
            n41367, n41441, n41229, n41227, n41319, w_result_sel_mul_d, 
            n41381, n41451, REF_CLK_c_enable_1030, n45106, REF_CLK_c_enable_1042, 
            REF_CLK_c_enable_1050, REF_CLK_c_enable_1299, \LM32I_ADR_O[4] , 
            \LM32I_ADR_O[5] , \LM32I_ADR_O[6] , \LM32I_ADR_O[7] , \LM32I_ADR_O[8] , 
            \LM32I_ADR_O[9] , \LM32I_ADR_O[10] , \LM32I_ADR_O[11] , \LM32I_ADR_O[12] , 
            \LM32I_ADR_O[13] , \LM32I_ADR_O[14] , \LM32I_ADR_O[15] , \LM32I_ADR_O[16] , 
            \LM32I_ADR_O[17] , \LM32I_ADR_O[18] , \LM32I_ADR_O[19] , \LM32I_ADR_O[20] , 
            \LM32I_ADR_O[21] , \LM32I_ADR_O[22] , \LM32I_ADR_O[23] , \LM32I_ADR_O[24] , 
            \LM32I_ADR_O[25] , \LM32I_ADR_O[26] , \LM32I_ADR_O[27] , \LM32I_ADR_O[28] , 
            \LM32I_ADR_O[29] , \LM32I_ADR_O[30] , \LM32I_ADR_O[31] , REF_CLK_c_enable_1425, 
            n41285, n30888, n41350, n41351, n41247, n41348, \instruction_d[11] , 
            \instruction_d[12] , \instruction_d[13] , \instruction_d[14] , 
            n41352, n41353, n41354, \write_idx_m[1] , n2_adj_166, 
            \write_idx_x[1] , n2_adj_167, n41355, n41356, n41357, 
            \write_idx_m[4] , n5, n41358, n45099, n2_adj_168, n41282, 
            n41359, n10475, n41366, n41368, n41369, n41370, n41371, 
            n41372, pc_a_31__N_1720, n41373, n41374, n41375, n41376, 
            n41377, n41179, \extended_immediate[31] , n2_adj_169, n41291, 
            n2_adj_170, n2_adj_171, n2_adj_172, n2_adj_173, n2_adj_174, 
            n2_adj_175, n2_adj_176, n6028, n41232, n35032, n12412, 
            dcache_refilling, dcache_refill_request, dcache_restart_request, 
            n949, n32220, locked_N_493, n40093, write_idx_d, n41380, 
            LM32D_CYC_O, n30879, n10485, n31519, selected, m_result_sel_shift_d, 
            n30058, n41362, LM32D_WE_O, \LM32D_ADR_O[1] , n41452, 
            n41241, n37918, n37916, n37917, n37919, n37915, n37914, 
            n36389, flush_set, icache_restart_request, restart_request_N_1998, 
            icache_refilling, \state[2] , n41196, n15, q_d, n45175, 
            valid_x_N_1285, n32278, n10_adj_177, n32264, n41203, n41408, 
            flush_set_8__N_1953, n9304, n41, n41187, branch_target_d, 
            n157, n31996, cycles_5__N_2934, REF_CLK_c_enable_1366, REF_CLK_c_enable_1622, 
            n41172, n32618, GND_net) /* synthesis syn_module_defined=1 */ ;
    output \genblk1.wait_one_tick_done ;
    output n6781;
    output n41208;
    output n6764;
    output n6769;
    output n6749;
    input REF_CLK_c;
    input stall_a;
    output way_match_0__N_2007;
    output bus_error_f_N_1884;
    output n41410;
    input n13990;
    input n32216;
    input n45075;
    input n41244;
    input n41419;
    output n41295;
    output n41248;
    output n30216;
    input REF_CLK_c_enable_1606;
    input VCC_net;
    input n41178;
    output \LM32I_CTI_O[0] ;
    input REF_CLK_c_enable_97;
    input n30900;
    output [31:2]pc_d;
    input REF_CLK_c_enable_1178;
    output [31:2]pc_f;
    output [31:2]pc_x;
    input REF_CLK_c_enable_1624;
    output [31:2]pc_m;
    input REF_CLK_c_enable_1235;
    input REF_CLK_c_enable_1131;
    input [31:0]SHAREDBUS_DAT_O;
    output n6760;
    output n6765;
    output n31717;
    output n45105;
    output n6771;
    input n73;
    output n41461;
    output n41228;
    output n41365;
    output n41361;
    output scall_d;
    output n41437;
    output n6778;
    output n6780;
    output n31542;
    output n6768;
    input n32910;
    output n6779;
    output n10;
    output n6777;
    output n6775;
    input branch_taken_m;
    output icache_refill_request;
    output \next_cycle_type[2] ;
    input n45080;
    input n41390;
    input n5223;
    output n37955;
    output n37956;
    output n37954;
    input n41345;
    output n41250;
    output n41251;
    output n41279;
    output \LM32I_ADR_O[2] ;
    input n45079;
    input \reg_12[2] ;
    output n2;
    input \reg_12[12] ;
    output n40677;
    input \reg_12[29] ;
    output n2_adj_149;
    input \reg_12[3] ;
    output n2_adj_150;
    input \reg_12[6] ;
    output n2_adj_151;
    input \reg_12[4] ;
    output n2_adj_152;
    input \reg_12[14] ;
    output n2_adj_153;
    input n30241;
    input n31750;
    input n31955;
    input n41429;
    input \reg_12[22] ;
    output n2_adj_154;
    input \reg_12[13] ;
    output n2_adj_155;
    input \reg_12[21] ;
    output n2_adj_156;
    input \reg_12[28] ;
    output n2_adj_157;
    input \reg_12[11] ;
    output n2_adj_158;
    input \reg_12[18] ;
    output n2_adj_159;
    input \reg_12[25] ;
    output n2_adj_160;
    input \reg_12[9] ;
    output n2_adj_161;
    input \reg_12[17] ;
    output n2_adj_162;
    input \reg_12[24] ;
    output n2_adj_163;
    input \reg_12[7] ;
    output n2_adj_164;
    input \reg_12[15] ;
    output n2_adj_165;
    output n41382;
    input n45183;
    output n6770;
    input n6589;
    input n6584;
    output n37179;
    input \write_idx_x[0] ;
    input n35751;
    output n35860;
    input n6439;
    input n6434;
    output n37177;
    input n6599;
    input n6594;
    output n37180;
    input n6629;
    input n6624;
    output n37183;
    input n6579;
    input n6574;
    output n37178;
    input n6429;
    input n6424;
    output n37176;
    input n45103;
    input n35687;
    output n35832;
    input n6609;
    input n6604;
    output n37181;
    input n6619;
    input n6614;
    output n37182;
    input n37185;
    input n37184;
    output n37188;
    input n37187;
    input n37186;
    output n37189;
    input n7603;
    input n7571;
    output [31:0]n7609;
    input n7607;
    input n7575;
    input n7606;
    input n7574;
    output bus_error_d;
    input n7604;
    input n7572;
    input n7605;
    input n7573;
    input n7608;
    input n7576;
    input n7602;
    input n7570;
    output \selected_1__N_354[0] ;
    input n7601;
    input n7569;
    input n7600;
    input n7568;
    input n7599;
    input n7567;
    input n7598;
    input n7566;
    input n7597;
    input n7565;
    input n7596;
    input n7564;
    input n7595;
    input n7563;
    input n7594;
    input n7562;
    input n7593;
    input n7561;
    input n7592;
    input n7560;
    input n7584;
    input n7552;
    input n7583;
    input n7551;
    input n7582;
    input n7550;
    input n7581;
    input n7549;
    input n7580;
    input n7548;
    input n7579;
    input n7547;
    input n7578;
    input n7546;
    input n7577;
    input n7545;
    output n6750;
    input n7591;
    input n7559;
    input n7590;
    input n7558;
    input n7589;
    input n7557;
    input n7588;
    input n7556;
    input n7587;
    input n7555;
    input n7586;
    input n7554;
    input n7585;
    input n7553;
    input n4;
    input \write_idx_x[3] ;
    output n32116;
    input n41430;
    input \write_idx_w[3] ;
    output n33920;
    output n37501;
    output n37500;
    output n37502;
    output n37499;
    output n37498;
    output n37497;
    output n37496;
    output n6751;
    output n6752;
    output n6753;
    output n6754;
    output n6755;
    output n6756;
    output n6757;
    output n6758;
    output n6759;
    output n6761;
    output n6762;
    output n6763;
    output n6766;
    output n6767;
    output n6776;
    input n40094;
    output n37495;
    input n7672;
    input n7640;
    output [31:0]n7677;
    input n7673;
    input n7641;
    input \write_idx_x[4] ;
    input n32260;
    output n32262;
    input n41312;
    output n41296;
    output n34;
    input n7674;
    input n7642;
    input n7675;
    input n7643;
    input n7676;
    input n7644;
    input n7671;
    input n7639;
    input n7670;
    input n7638;
    input n7669;
    input n7637;
    input n7668;
    input n7636;
    input n7667;
    input n7635;
    input n7666;
    input n7634;
    input n7665;
    input n7633;
    input n7664;
    input n7632;
    input n7663;
    input n7631;
    input n7662;
    input n7630;
    input n7661;
    input n7629;
    input n7660;
    input n7628;
    output n36;
    input n7652;
    input n7620;
    input n7651;
    input n7619;
    input n7650;
    input n7618;
    input n7649;
    input n7617;
    output n37;
    input n7648;
    input n7616;
    input n7647;
    input n7615;
    input n7646;
    input n7614;
    input n7645;
    input n7613;
    input n7659;
    input n7627;
    input n7658;
    input n7626;
    input n7657;
    input n7625;
    input n7656;
    input n7624;
    input n7655;
    input n7623;
    input n7654;
    input n7622;
    input n7653;
    input n7621;
    input n30012;
    input \write_idx_m[2] ;
    output n31976;
    input n37504;
    input n37503;
    output n37507;
    input n37506;
    input n37505;
    output n37508;
    input n41364;
    output n41363;
    output n30820;
    input n11834;
    output n41216;
    input n32356;
    output n41281;
    output n41367;
    input n41441;
    output n41229;
    output n41227;
    input n41319;
    output w_result_sel_mul_d;
    output n41381;
    input n41451;
    input REF_CLK_c_enable_1030;
    output n45106;
    input REF_CLK_c_enable_1042;
    input REF_CLK_c_enable_1050;
    input REF_CLK_c_enable_1299;
    output \LM32I_ADR_O[4] ;
    output \LM32I_ADR_O[5] ;
    output \LM32I_ADR_O[6] ;
    output \LM32I_ADR_O[7] ;
    output \LM32I_ADR_O[8] ;
    output \LM32I_ADR_O[9] ;
    output \LM32I_ADR_O[10] ;
    output \LM32I_ADR_O[11] ;
    output \LM32I_ADR_O[12] ;
    output \LM32I_ADR_O[13] ;
    output \LM32I_ADR_O[14] ;
    output \LM32I_ADR_O[15] ;
    output \LM32I_ADR_O[16] ;
    output \LM32I_ADR_O[17] ;
    output \LM32I_ADR_O[18] ;
    output \LM32I_ADR_O[19] ;
    output \LM32I_ADR_O[20] ;
    output \LM32I_ADR_O[21] ;
    output \LM32I_ADR_O[22] ;
    output \LM32I_ADR_O[23] ;
    output \LM32I_ADR_O[24] ;
    output \LM32I_ADR_O[25] ;
    output \LM32I_ADR_O[26] ;
    output \LM32I_ADR_O[27] ;
    output \LM32I_ADR_O[28] ;
    output \LM32I_ADR_O[29] ;
    output \LM32I_ADR_O[30] ;
    output \LM32I_ADR_O[31] ;
    input REF_CLK_c_enable_1425;
    output n41285;
    output n30888;
    output n41350;
    output n41351;
    output n41247;
    output n41348;
    output \instruction_d[11] ;
    output \instruction_d[12] ;
    output \instruction_d[13] ;
    output \instruction_d[14] ;
    output n41352;
    output n41353;
    output n41354;
    input \write_idx_m[1] ;
    output n2_adj_166;
    input \write_idx_x[1] ;
    output n2_adj_167;
    output n41355;
    output n41356;
    output n41357;
    input \write_idx_m[4] ;
    output n5;
    output n41358;
    input n45099;
    output n2_adj_168;
    output n41282;
    output n41359;
    input n10475;
    output n41366;
    output n41368;
    output n41369;
    output n41370;
    output n41371;
    output n41372;
    input [29:0]pc_a_31__N_1720;
    output n41373;
    output n41374;
    output n41375;
    output n41376;
    output n41377;
    input n41179;
    input \extended_immediate[31] ;
    input n2_adj_169;
    input n41291;
    output n2_adj_170;
    input n2_adj_171;
    output n2_adj_172;
    input n2_adj_173;
    output n2_adj_174;
    input n2_adj_175;
    output n2_adj_176;
    output n6028;
    input n41232;
    input n35032;
    output n12412;
    input dcache_refilling;
    input dcache_refill_request;
    input dcache_restart_request;
    input [0:0]n949;
    input n32220;
    output locked_N_493;
    output n40093;
    output [4:0]write_idx_d;
    input n41380;
    input LM32D_CYC_O;
    output n30879;
    input n10485;
    output n31519;
    input [1:0]selected;
    output m_result_sel_shift_d;
    input n30058;
    output n41362;
    input LM32D_WE_O;
    input \LM32D_ADR_O[1] ;
    output n41452;
    output n41241;
    input n37918;
    input n37916;
    input n37917;
    input n37919;
    input n37915;
    input n37914;
    input n36389;
    output [8:0]flush_set;
    output icache_restart_request;
    input restart_request_N_1998;
    output icache_refilling;
    output \state[2] ;
    input n41196;
    input n15;
    input q_d;
    input n45175;
    output valid_x_N_1285;
    input n32278;
    input n10_adj_177;
    input n32264;
    input n41203;
    input n41408;
    input [8:0]flush_set_8__N_1953;
    output n9304;
    output n41;
    input n41187;
    input [31:2]branch_target_d;
    input [29:0]n157;
    input n31996;
    input cycles_5__N_2934;
    output REF_CLK_c_enable_1366;
    output REF_CLK_c_enable_1622;
    input n41172;
    input n32618;
    input GND_net;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    
    wire n41475, n41474, n40272, n12048, n20031, n29933;
    wire [29:0]pc_a_31__N_1598;
    wire [31:2]restart_address;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(337[20:35])
    wire [31:2]pc_a;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(334[20:24])
    wire [31:2]pc_w;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(260[23:27])
    
    wire REF_CLK_c_enable_1100;
    wire [29:0]restart_address_31__N_1628;
    wire [31:0]icache_refill_data;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(344[29:47])
    
    wire bus_error_f, REF_CLK_c_enable_129, n41478, n41477, n32670, 
        n6772, n6773, n6774, n41459, n41460, n32152, n7077, n7045;
    wire [10:0]\genblk1.ra ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(285[31:33])
    
    wire n40069, n41471, n32046, icache_refill_ready, n38967, n38966, 
        n7155, n7123, n40068, n40179, n40180, n40149, n40150, 
        n40136, n40137, n40126, n40127, REF_CLK_c_enable_406, n9336, 
        n7156, n7124, n40073, n7078, n7046, n40074, n40233, n40131, 
        n40132, n40141, n40142, n40174, n40175, n7143, n7175, 
        n40091, n7065, n7097, n40090, n40228, n40223, n40215, 
        n40210, n40205, n40200, n40195, n40190, n40185, n40072, 
        n40077, n40238, n40281, n40170, n40165, n40160, n40155, 
        n40122, n40117, n40112, n40107, n40099, n7064, n7096, 
        n40095, n40159, n7142, n7174, n40096, n40154, n7141, n7173, 
        n40104, n7063, n7095, n40103, n7062, n7094, n40108, n7140, 
        n7172, n40109, n40169, n7061, n7093, n40113, n40164, n7139, 
        n7171, n40114, n7060, n7092, n40118, n7138, n7170, n40119, 
        n40227, n40280, n45201, n40098, n7059, n7091, n40123, 
        n7137, n7169, n40124, n7058, n7090, n40128, n40106, n7136, 
        n7168, n40129, n7057, n7089, n40133, n7135, n7167, n40134, 
        n40121, n7056, n7088, n40138, n7134, n7166, n40139, n40116, 
        n7133, n7165, n40147, n7055, n7087, n40146, n7054, n7086, 
        n40151, n7132, n7164, n40152, n40278, n40277, n40279, 
        n40270, n40268, n37144, n40271, n7053, n7085, n40156, 
        n7131, n7163, n40157, n40232, n40222, n7052, n7084, n40161, 
        n40214, n40209, n7130, n7162, n40162, n40204, n40199, 
        n40194, n40189, n40184, n40237, n45202, n7051, n7083, 
        n40166, n7129, n7161, n40167, n7050, n7082, n40171, n40235, 
        n40234, n40236, n7128, n7160, n40172, n7049, n7081, n40176, 
        n7127, n7159, n40177, n7044, n7076, n40181, n7122, n7154, 
        n40182, REF_CLK_c_enable_1133;
    wire [31:0]i_adr_o_31__N_1531;
    
    wire n40231, n40229, n7043, n7075, n40186, n40226, n40224, 
        REF_CLK_c_enable_1161;
    wire [31:2]icache_refill_address;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(342[21:42])
    
    wire n7121, n7153, n40187, n40221, n40219, n40213, n40211, 
        n7042, n7074, n40191, n7120, n7152, n40192, n40208, n40206, 
        n7041, n7073, n40196, n40203, n40201, n45204, n45205, 
        n7119, n7151, n40197, n40198, n7040, n7072, n7118, n7150, 
        n40202, n7039, n7071, n41465, n40193, n7117, n7149, n40207, 
        n40188, n7038, n7070, n7116, n7148, n40212, n40183, n40178, 
        n7115, n7147, n40220, n7037, n7069, n40173, n40168, n40163, 
        n7036, n7068, n40158, n7114, n7146, n40225, n40153, n40148, 
        n40140, n7035, n7067, n7113, n7145, n40230, n40135, n7157, 
        n7125, n7079, n7047, n40130, n40125, n40120, n40115, n40110, 
        n40111, n31807, n35314, n7112, n7144, n40269, n41469, 
        n40105, n41468, n7034, n7066, n40097, n40092, n7080, n7048, 
        n40076, n40075, n7158, n7126, n40071, n41472, n40070, 
        n32478;
    wire [29:0]pc_a_31__N_1690;
    
    wire n41466, n1;
    
    LUT4 i15103_3_lut_4_lut_then_4_lut (.A(\genblk1.wait_one_tick_done ), 
         .B(n6781), .C(n41208), .D(n6764), .Z(n41475)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i15103_3_lut_4_lut_then_4_lut.init = 16'h2f0f;
    LUT4 i15103_3_lut_4_lut_else_4_lut (.A(\genblk1.wait_one_tick_done ), 
         .B(n6781), .C(n41208), .D(n6769), .Z(n41474)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i15103_3_lut_4_lut_else_4_lut.init = 16'h2f0f;
    FD1S3AX instruction_d__2828_rep_4_i1 (.D(n40272), .CK(REF_CLK_c), .Q(n6749)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i1.GSR = "ENABLED";
    FD1S3IX instruction_d__2828 (.D(way_match_0__N_2007), .CK(REF_CLK_c), 
            .CD(stall_a), .Q(n6781));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828.GSR = "ENABLED";
    LUT4 i1_4_lut_4_lut (.A(bus_error_f_N_1884), .B(n41410), .C(n13990), 
         .D(n32216), .Z(n12048)) /* synthesis lut_function=(A ((D)+!C)+!A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i1_4_lut_4_lut.init = 16'hee4e;
    LUT4 i1_4_lut (.A(n45075), .B(n41244), .C(n20031), .D(n41419), .Z(n29933)) /* synthesis lut_function=(A (B+(D))+!A !(B (C)+!B (C+!(D)))) */ ;
    defparam i1_4_lut.init = 16'haf8c;
    LUT4 i25200_4_lut (.A(n41295), .B(n20031), .C(n41248), .D(n41244), 
         .Z(n30216)) /* synthesis lut_function=(A (B)+!A (B+!(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(460[6:19])
    defparam i25200_4_lut.init = 16'hcddd;
    FD1S3DX \genblk1.wait_one_tick_done_270  (.D(VCC_net), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\genblk1.wait_one_tick_done )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(418[12] 423[38])
    defparam \genblk1.wait_one_tick_done_270 .GSR = "ENABLED";
    LUT4 pc_a_31__I_0_i6_rep_123_3_lut (.A(pc_a_31__N_1598[5]), .B(restart_address[7]), 
         .C(n41178), .Z(pc_a[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(493[7] 511[25])
    defparam pc_a_31__I_0_i6_rep_123_3_lut.init = 16'hcaca;
    FD1P3BX i_cti_o__i1 (.D(n30900), .SP(REF_CLK_c_enable_97), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(\LM32I_CTI_O[0] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_cti_o__i1.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i2 (.D(pc_f[2]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i2.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i2 (.D(pc_d[2]), .SP(REF_CLK_c_enable_1624), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i2.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i2 (.D(pc_x[2]), .SP(REF_CLK_c_enable_1235), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i2.GSR = "ENABLED";
    FD1S3DX pc_w_i2 (.D(pc_m[2]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i2.GSR = "ENABLED";
    FD1P3DX restart_address_i2 (.D(restart_address_31__N_1628[0]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i2.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i0 (.D(SHAREDBUS_DAT_O[0]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i0.GSR = "ENABLED";
    FD1P3BX pc_f_i2_i2 (.D(pc_a[2]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(pc_f[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i2.GSR = "ENABLED";
    FD1P3DX bus_error_f_116 (.D(bus_error_f_N_1884), .SP(REF_CLK_c_enable_129), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(bus_error_f)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam bus_error_f_116.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut_then_4_lut (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n41208), .D(n6760), .Z(n41478)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_3_lut_4_lut_then_4_lut.init = 16'h2f0f;
    LUT4 i1_3_lut_4_lut_else_4_lut (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n41208), .D(n6765), .Z(n41477)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_3_lut_4_lut_else_4_lut.init = 16'h2f0f;
    LUT4 i1_4_lut_adj_374 (.A(n32670), .B(n6781), .C(n6772), .D(n6773), 
         .Z(n31717)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(418[12] 423[38])
    defparam i1_4_lut_adj_374.init = 16'h2000;
    LUT4 i1_3_lut (.A(n6774), .B(n45105), .C(n6771), .Z(n32670)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(418[12] 423[38])
    defparam i1_3_lut.init = 16'h8080;
    PFUMX i34359 (.BLUT(n41459), .ALUT(n41460), .C0(n73), .Z(n41461));
    LUT4 i1_4_lut_adj_375 (.A(n32152), .B(n41228), .C(n41365), .D(n41361), 
         .Z(scall_d)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_4_lut_adj_375.init = 16'h2000;
    LUT4 n7077_bdd_3_lut (.A(n7077), .B(n7045), .C(\genblk1.ra [9]), .Z(n40069)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n7077_bdd_3_lut.init = 16'hacac;
    LUT4 i1_4_lut_adj_376 (.A(n41437), .B(n6781), .C(n6778), .D(n6780), 
         .Z(n31542)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_4_lut_adj_376.init = 16'h2000;
    LUT4 i1_3_lut_4_lut_else_4_lut_adj_377 (.A(\genblk1.wait_one_tick_done ), 
         .B(n6781), .C(n41208), .D(n6768), .Z(n41471)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_3_lut_4_lut_else_4_lut_adj_377.init = 16'h2f0f;
    LUT4 i1_4_lut_adj_378 (.A(n32910), .B(n6781), .C(n45105), .D(n6779), 
         .Z(n10)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_4_lut_adj_378.init = 16'h3020;
    LUT4 i1_2_lut (.A(n6777), .B(n6775), .Z(n32046)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 bus_error_f_N_1884_bdd_3_lut (.A(branch_taken_m), .B(icache_refill_ready), 
         .C(icache_refill_request), .Z(n38967)) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam bus_error_f_N_1884_bdd_3_lut.init = 16'hbaba;
    FD1S3DX icache_refill_ready_115 (.D(REF_CLK_c_enable_1131), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(icache_refill_ready)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_ready_115.GSR = "ENABLED";
    LUT4 i33195_rep_191_2_lut_4_lut (.A(\next_cycle_type[2] ), .B(n45080), 
         .C(n41390), .D(n5223), .Z(n37955)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i33195_rep_191_2_lut_4_lut.init = 16'hffca;
    LUT4 i33195_rep_192_2_lut_4_lut (.A(\next_cycle_type[2] ), .B(n45080), 
         .C(n41390), .D(n5223), .Z(n37956)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i33195_rep_192_2_lut_4_lut.init = 16'hffca;
    LUT4 i33195_rep_190_2_lut_4_lut (.A(\next_cycle_type[2] ), .B(n45080), 
         .C(n41390), .D(n5223), .Z(n37954)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i33195_rep_190_2_lut_4_lut.init = 16'hffca;
    LUT4 SPI_ADR_I_7__I_0_314_i10_2_lut_rep_845_4_lut (.A(\next_cycle_type[2] ), 
         .B(n45080), .C(n41390), .D(n41345), .Z(n41250)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B)) */ ;
    defparam SPI_ADR_I_7__I_0_314_i10_2_lut_rep_845_4_lut.init = 16'hff35;
    LUT4 SPI_ADR_I_7__I_0_313_i10_2_lut_rep_846_4_lut (.A(\next_cycle_type[2] ), 
         .B(n45080), .C(n41390), .D(n41345), .Z(n41251)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;
    defparam SPI_ADR_I_7__I_0_313_i10_2_lut_rep_846_4_lut.init = 16'hcaff;
    LUT4 equal_19_i3_2_lut_rep_874_4_lut (.A(\next_cycle_type[2] ), .B(n45080), 
         .C(n41390), .D(n41345), .Z(n41279)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam equal_19_i3_2_lut_rep_874_4_lut.init = 16'hffca;
    LUT4 i15227_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[2] ), .Z(n2)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15227_2_lut_4_lut.init = 16'hca00;
    LUT4 SHAREDBUS_ADR_I_3__bdd_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), 
         .C(n41390), .D(\reg_12[12] ), .Z(n40677)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam SHAREDBUS_ADR_I_3__bdd_2_lut_4_lut.init = 16'hca00;
    LUT4 i15200_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[29] ), .Z(n2_adj_149)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15200_2_lut_4_lut.init = 16'hca00;
    LUT4 i15226_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[3] ), .Z(n2_adj_150)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15226_2_lut_4_lut.init = 16'hca00;
    LUT4 i15223_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[6] ), .Z(n2_adj_151)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15223_2_lut_4_lut.init = 16'hca00;
    LUT4 i15225_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[4] ), .Z(n2_adj_152)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15225_2_lut_4_lut.init = 16'hca00;
    LUT4 i15215_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[14] ), .Z(n2_adj_153)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15215_2_lut_4_lut.init = 16'hca00;
    LUT4 bus_error_f_N_1884_bdd_4_lut (.A(n30241), .B(n31750), .C(n31955), 
         .D(n41429), .Z(n38966)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam bus_error_f_N_1884_bdd_4_lut.init = 16'h0200;
    LUT4 i15207_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[22] ), .Z(n2_adj_154)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15207_2_lut_4_lut.init = 16'hca00;
    LUT4 i15216_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[13] ), .Z(n2_adj_155)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15216_2_lut_4_lut.init = 16'hca00;
    LUT4 i15208_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[21] ), .Z(n2_adj_156)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15208_2_lut_4_lut.init = 16'hca00;
    LUT4 i15201_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[28] ), .Z(n2_adj_157)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15201_2_lut_4_lut.init = 16'hca00;
    LUT4 i15218_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[11] ), .Z(n2_adj_158)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15218_2_lut_4_lut.init = 16'hca00;
    LUT4 i15211_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[18] ), .Z(n2_adj_159)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15211_2_lut_4_lut.init = 16'hca00;
    LUT4 i15204_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[25] ), .Z(n2_adj_160)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15204_2_lut_4_lut.init = 16'hca00;
    LUT4 i15220_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[9] ), .Z(n2_adj_161)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15220_2_lut_4_lut.init = 16'hca00;
    LUT4 i15212_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[17] ), .Z(n2_adj_162)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15212_2_lut_4_lut.init = 16'hca00;
    LUT4 i15205_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[24] ), .Z(n2_adj_163)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15205_2_lut_4_lut.init = 16'hca00;
    LUT4 i15222_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[7] ), .Z(n2_adj_164)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15222_2_lut_4_lut.init = 16'hca00;
    LUT4 n7077_bdd_3_lut_33948 (.A(n7155), .B(n7123), .C(\genblk1.ra [9]), 
         .Z(n40068)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n7077_bdd_3_lut_33948.init = 16'hacac;
    LUT4 i15214_2_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(n45079), .C(n41390), 
         .D(\reg_12[15] ), .Z(n2_adj_165)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i15214_2_lut_4_lut.init = 16'hca00;
    LUT4 n40179_bdd_3_lut_4_lut (.A(n41382), .B(n6764), .C(n45183), .D(n40179), 
         .Z(n40180)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40179_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n40149_bdd_3_lut_4_lut (.A(n6770), .B(n41382), .C(n45183), .D(n40149), 
         .Z(n40150)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40149_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i32007_3_lut_4_lut (.A(n6770), .B(n41382), .C(n6589), .D(n6584), 
         .Z(n37179)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32007_3_lut_4_lut.init = 16'hf780;
    LUT4 i30698_3_lut_4_lut (.A(n6770), .B(n41382), .C(\write_idx_x[0] ), 
         .D(n35751), .Z(n35860)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+(D)))+!A (C+(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i30698_3_lut_4_lut.init = 16'hff78;
    LUT4 i32005_3_lut_4_lut (.A(n6770), .B(n41382), .C(n6439), .D(n6434), 
         .Z(n37177)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32005_3_lut_4_lut.init = 16'hf780;
    LUT4 i32008_3_lut_4_lut (.A(n6770), .B(n41382), .C(n6599), .D(n6594), 
         .Z(n37180)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32008_3_lut_4_lut.init = 16'hf780;
    LUT4 i32011_3_lut_4_lut (.A(n6770), .B(n41382), .C(n6629), .D(n6624), 
         .Z(n37183)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32011_3_lut_4_lut.init = 16'hf780;
    LUT4 i32006_3_lut_4_lut (.A(n6770), .B(n41382), .C(n6579), .D(n6574), 
         .Z(n37178)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32006_3_lut_4_lut.init = 16'hf780;
    LUT4 i32004_3_lut_4_lut (.A(n6770), .B(n41382), .C(n6429), .D(n6424), 
         .Z(n37176)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32004_3_lut_4_lut.init = 16'hf780;
    LUT4 i30670_3_lut_4_lut (.A(n6770), .B(n41382), .C(n45103), .D(n35687), 
         .Z(n35832)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+(D)))+!A (C+(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i30670_3_lut_4_lut.init = 16'hff78;
    LUT4 i32009_3_lut_4_lut (.A(n6770), .B(n41382), .C(n6609), .D(n6604), 
         .Z(n37181)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32009_3_lut_4_lut.init = 16'hf780;
    LUT4 i32010_3_lut_4_lut (.A(n6770), .B(n41382), .C(n6619), .D(n6614), 
         .Z(n37182)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32010_3_lut_4_lut.init = 16'hf780;
    LUT4 n40136_bdd_3_lut_4_lut (.A(n41382), .B(n6772), .C(n45183), .D(n40136), 
         .Z(n40137)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n40136_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i32016_3_lut_4_lut (.A(n41382), .B(n6772), .C(n37185), .D(n37184), 
         .Z(n37188)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i32016_3_lut_4_lut.init = 16'hf780;
    LUT4 i32017_3_lut_4_lut (.A(n41382), .B(n6772), .C(n37187), .D(n37186), 
         .Z(n37189)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i32017_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i27_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7603), .D(n7571), 
         .Z(n7609[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i27_3_lut_4_lut.init = 16'hf780;
    LUT4 n40126_bdd_3_lut_4_lut (.A(n41382), .B(n6774), .C(n45183), .D(n40126), 
         .Z(n40127)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n40126_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_3145_i31_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7607), .D(n7575), 
         .Z(n7609[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i31_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i30_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7606), .D(n7574), 
         .Z(n7609[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i30_3_lut_4_lut.init = 16'hf780;
    FD1P3DX bus_error_d_118 (.D(bus_error_f), .SP(REF_CLK_c_enable_1178), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(bus_error_d)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam bus_error_d_118.GSR = "ENABLED";
    FD1S3DX i_cyc_o_109 (.D(n12048), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(bus_error_f_N_1884)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_cyc_o_109.GSR = "ENABLED";
    LUT4 mux_3145_i28_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7604), .D(n7572), 
         .Z(n7609[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i28_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i29_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7605), .D(n7573), 
         .Z(n7609[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i29_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i32_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7608), .D(n7576), 
         .Z(n7609[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i32_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i26_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7602), .D(n7570), 
         .Z(n7609[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i26_3_lut_4_lut.init = 16'hf780;
    FD1P3DX i_stb_o_110 (.D(n9336), .SP(REF_CLK_c_enable_406), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\selected_1__N_354[0] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_stb_o_110.GSR = "ENABLED";
    LUT4 mux_3145_i25_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7601), .D(n7569), 
         .Z(n7609[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i25_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i24_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7600), .D(n7568), 
         .Z(n7609[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i24_3_lut_4_lut.init = 16'hf780;
    LUT4 pc_a_31__I_0_i8_rep_131_3_lut (.A(pc_a_31__N_1598[7]), .B(restart_address[9]), 
         .C(n41178), .Z(pc_a[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(493[7] 511[25])
    defparam pc_a_31__I_0_i8_rep_131_3_lut.init = 16'hcaca;
    LUT4 mux_3145_i23_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7599), .D(n7567), 
         .Z(n7609[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i23_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i22_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7598), .D(n7566), 
         .Z(n7609[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i21_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7597), .D(n7565), 
         .Z(n7609[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i20_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7596), .D(n7564), 
         .Z(n7609[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i19_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7595), .D(n7563), 
         .Z(n7609[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i18_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7594), .D(n7562), 
         .Z(n7609[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i17_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7593), .D(n7561), 
         .Z(n7609[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i16_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7592), .D(n7560), 
         .Z(n7609[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i8_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7584), .D(n7552), 
         .Z(n7609[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i7_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7583), .D(n7551), 
         .Z(n7609[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 n7078_bdd_3_lut_33953 (.A(n7156), .B(n7124), .C(\genblk1.ra [9]), 
         .Z(n40073)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n7078_bdd_3_lut_33953.init = 16'hacac;
    LUT4 mux_3145_i6_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7582), .D(n7550), 
         .Z(n7609[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 n7078_bdd_3_lut (.A(n7078), .B(n7046), .C(\genblk1.ra [9]), .Z(n40074)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n7078_bdd_3_lut.init = 16'hacac;
    LUT4 mux_3145_i5_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7581), .D(n7549), 
         .Z(n7609[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i4_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7580), .D(n7548), 
         .Z(n7609[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i3_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7579), .D(n7547), 
         .Z(n7609[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i2_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7578), .D(n7546), 
         .Z(n7609[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i1_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7577), .D(n7545), 
         .Z(n7609[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i1_3_lut_4_lut.init = 16'hf780;
    FD1S3AX instruction_d__2828_rep_4_i2 (.D(n40233), .CK(REF_CLK_c), .Q(n6750)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i2.GSR = "ENABLED";
    LUT4 mux_3145_i15_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7591), .D(n7559), 
         .Z(n7609[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i14_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7590), .D(n7558), 
         .Z(n7609[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i13_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7589), .D(n7557), 
         .Z(n7609[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i12_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7588), .D(n7556), 
         .Z(n7609[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i11_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7587), .D(n7555), 
         .Z(n7609[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i10_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7586), .D(n7554), 
         .Z(n7609[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3145_i9_3_lut_4_lut (.A(n41382), .B(n6774), .C(n7585), .D(n7553), 
         .Z(n7609[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_3145_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 n40131_bdd_3_lut_4_lut (.A(n41382), .B(n6773), .C(n45183), .D(n40131), 
         .Z(n40132)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n40131_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_3_lut_4_lut (.A(n41382), .B(n6773), .C(n4), .D(\write_idx_x[3] ), 
         .Z(n32116)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h8070;
    LUT4 i1_3_lut_4_lut_adj_379 (.A(n41382), .B(n6773), .C(n41430), .D(\write_idx_w[3] ), 
         .Z(n33920)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam i1_3_lut_4_lut_adj_379.init = 16'h8070;
    LUT4 n40141_bdd_3_lut_4_lut (.A(n6771), .B(n41382), .C(n45183), .D(n40141), 
         .Z(n40142)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40141_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n40174_bdd_3_lut_4_lut (.A(n6765), .B(n41382), .C(n45183), .D(n40174), 
         .Z(n40175)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40174_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i32329_3_lut_4_lut (.A(n6765), .B(n41382), .C(n6619), .D(n6614), 
         .Z(n37501)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32329_3_lut_4_lut.init = 16'hf780;
    LUT4 i32328_3_lut_4_lut (.A(n6765), .B(n41382), .C(n6609), .D(n6604), 
         .Z(n37500)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32328_3_lut_4_lut.init = 16'hf780;
    LUT4 n6874_bdd_3_lut_33961 (.A(n7143), .B(\genblk1.ra [9]), .C(n7175), 
         .Z(n40091)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33961.init = 16'he2e2;
    LUT4 i32330_3_lut_4_lut (.A(n6765), .B(n41382), .C(n6629), .D(n6624), 
         .Z(n37502)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32330_3_lut_4_lut.init = 16'hf780;
    LUT4 i32327_3_lut_4_lut (.A(n6765), .B(n41382), .C(n6599), .D(n6594), 
         .Z(n37499)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32327_3_lut_4_lut.init = 16'hf780;
    LUT4 i32326_3_lut_4_lut (.A(n6765), .B(n41382), .C(n6589), .D(n6584), 
         .Z(n37498)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32326_3_lut_4_lut.init = 16'hf780;
    LUT4 i32325_3_lut_4_lut (.A(n6765), .B(n41382), .C(n6579), .D(n6574), 
         .Z(n37497)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32325_3_lut_4_lut.init = 16'hf780;
    LUT4 i32324_3_lut_4_lut (.A(n6765), .B(n41382), .C(n6439), .D(n6434), 
         .Z(n37496)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32324_3_lut_4_lut.init = 16'hf780;
    LUT4 n6874_bdd_3_lut_33958 (.A(n7065), .B(\genblk1.ra [9]), .C(n7097), 
         .Z(n40090)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33958.init = 16'he2e2;
    FD1S3AX instruction_d__2828_rep_4_i3 (.D(n40228), .CK(REF_CLK_c), .Q(n6751)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i3.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i4 (.D(n40223), .CK(REF_CLK_c), .Q(n6752)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i4.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i5 (.D(n40215), .CK(REF_CLK_c), .Q(n6753)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i5.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i6 (.D(n40210), .CK(REF_CLK_c), .Q(n6754)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i6.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i7 (.D(n40205), .CK(REF_CLK_c), .Q(n6755)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i7.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i8 (.D(n40200), .CK(REF_CLK_c), .Q(n6756)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i8.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i9 (.D(n40195), .CK(REF_CLK_c), .Q(n6757)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i9.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i10 (.D(n40190), .CK(REF_CLK_c), .Q(n6758)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i10.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i11 (.D(n40185), .CK(REF_CLK_c), .Q(n6759)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i11.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i12 (.D(n40072), .CK(REF_CLK_c), .Q(n6760)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i12.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i13 (.D(n40077), .CK(REF_CLK_c), .Q(n6761)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i13.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i14 (.D(n40238), .CK(REF_CLK_c), .Q(n6762)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i14.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i15 (.D(n40281), .CK(REF_CLK_c), .Q(n6763)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i15.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i16 (.D(n40180), .CK(REF_CLK_c), .Q(n6764)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i16.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i17 (.D(n40175), .CK(REF_CLK_c), .Q(n6765)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i17.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i18 (.D(n40170), .CK(REF_CLK_c), .Q(n6766)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i18.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i19 (.D(n40165), .CK(REF_CLK_c), .Q(n6767)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i19.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i20 (.D(n40160), .CK(REF_CLK_c), .Q(n6768)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i20.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i21 (.D(n40155), .CK(REF_CLK_c), .Q(n6769)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i21.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i22 (.D(n40150), .CK(REF_CLK_c), .Q(n6770)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i22.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i23 (.D(n40142), .CK(REF_CLK_c), .Q(n6771)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i23.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i24 (.D(n40137), .CK(REF_CLK_c), .Q(n6772)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i24.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i25 (.D(n40132), .CK(REF_CLK_c), .Q(n6773)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i25.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i26 (.D(n40127), .CK(REF_CLK_c), .Q(n6774)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i26.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i27 (.D(n40122), .CK(REF_CLK_c), .Q(n6775)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i27.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i28 (.D(n40117), .CK(REF_CLK_c), .Q(n6776)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i28.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i29 (.D(n40112), .CK(REF_CLK_c), .Q(n6777)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i29.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i30 (.D(n40107), .CK(REF_CLK_c), .Q(n6778)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i30.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i31 (.D(n40099), .CK(REF_CLK_c), .Q(n6779)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i31.GSR = "ENABLED";
    FD1S3AX instruction_d__2828_rep_4_i32 (.D(n40094), .CK(REF_CLK_c), .Q(n6780)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d__2828_rep_4_i32.GSR = "ENABLED";
    LUT4 i32323_3_lut_4_lut (.A(n6765), .B(n41382), .C(n6429), .D(n6424), 
         .Z(n37495)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32323_3_lut_4_lut.init = 16'hf780;
    LUT4 pc_a_31__I_0_i7_rep_127_3_lut (.A(pc_a_31__N_1598[6]), .B(restart_address[8]), 
         .C(n41178), .Z(pc_a[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(493[7] 511[25])
    defparam pc_a_31__I_0_i7_rep_127_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_0_i5_rep_129_3_lut (.A(pc_a_31__N_1598[4]), .B(restart_address[6]), 
         .C(n41178), .Z(pc_a[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(493[7] 511[25])
    defparam pc_a_31__I_0_i5_rep_129_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_0_i3_rep_125_3_lut (.A(pc_a_31__N_1598[2]), .B(restart_address[4]), 
         .C(n41178), .Z(pc_a[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(493[7] 511[25])
    defparam pc_a_31__I_0_i3_rep_125_3_lut.init = 16'hcaca;
    LUT4 n6874_bdd_3_lut_33962 (.A(n7064), .B(\genblk1.ra [9]), .C(n7096), 
         .Z(n40095)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33962.init = 16'he2e2;
    LUT4 n40159_bdd_3_lut_4_lut (.A(n6768), .B(n41382), .C(n45183), .D(n40159), 
         .Z(n40160)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40159_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n6874_bdd_3_lut_33965 (.A(n7142), .B(\genblk1.ra [9]), .C(n7174), 
         .Z(n40096)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33965.init = 16'he2e2;
    LUT4 mux_3183_i28_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7672), .D(n7640), 
         .Z(n7677[27])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i28_3_lut_4_lut.init = 16'hf780;
    LUT4 n40154_bdd_3_lut_4_lut (.A(n6769), .B(n41382), .C(n45183), .D(n40154), 
         .Z(n40155)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40154_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_3183_i29_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7673), .D(n7641), 
         .Z(n7677[28])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i29_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_3_lut_4_lut_adj_380 (.A(n6769), .B(n41382), .C(\write_idx_x[4] ), 
         .D(n32260), .Z(n32262)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+(D)))+!A (C+(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_3_lut_4_lut_adj_380.init = 16'hff78;
    LUT4 i1_3_lut_4_lut_adj_381 (.A(n41312), .B(n6764), .C(n6774), .D(n41296), 
         .Z(n34)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_3_lut_4_lut_adj_381.init = 16'hf888;
    LUT4 mux_3183_i30_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7674), .D(n7642), 
         .Z(n7677[29])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i30_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i31_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7675), .D(n7643), 
         .Z(n7677[30])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i31_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i32_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7676), .D(n7644), 
         .Z(n7677[31])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i32_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i27_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7671), .D(n7639), 
         .Z(n7677[26])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i27_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i26_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7670), .D(n7638), 
         .Z(n7677[25])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i26_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i25_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7669), .D(n7637), 
         .Z(n7677[24])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i25_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i24_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7668), .D(n7636), 
         .Z(n7677[23])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i24_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i23_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7667), .D(n7635), 
         .Z(n7677[22])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i23_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i22_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7666), .D(n7634), 
         .Z(n7677[21])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 n6874_bdd_3_lut_33969 (.A(n7141), .B(\genblk1.ra [9]), .C(n7173), 
         .Z(n40104)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33969.init = 16'he2e2;
    LUT4 mux_3183_i21_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7665), .D(n7633), 
         .Z(n7677[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 n6874_bdd_3_lut_33966 (.A(n7063), .B(\genblk1.ra [9]), .C(n7095), 
         .Z(n40103)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33966.init = 16'he2e2;
    LUT4 mux_3183_i20_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7664), .D(n7632), 
         .Z(n7677[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i19_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7663), .D(n7631), 
         .Z(n7677[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i18_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7662), .D(n7630), 
         .Z(n7677[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i17_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7661), .D(n7629), 
         .Z(n7677[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i16_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7660), .D(n7628), 
         .Z(n7677[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_3_lut_4_lut_adj_382 (.A(n41312), .B(n6764), .C(n6772), .D(n41296), 
         .Z(n36)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_3_lut_4_lut_adj_382.init = 16'hf888;
    LUT4 mux_3183_i8_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7652), .D(n7620), 
         .Z(n7677[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i7_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7651), .D(n7619), 
         .Z(n7677[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i6_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7650), .D(n7618), 
         .Z(n7677[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i5_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7649), .D(n7617), 
         .Z(n7677[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_3_lut_4_lut_adj_383 (.A(n41312), .B(n6764), .C(n6773), .D(n41296), 
         .Z(n37)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_3_lut_4_lut_adj_383.init = 16'hf888;
    LUT4 mux_3183_i4_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7648), .D(n7616), 
         .Z(n7677[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i3_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7647), .D(n7615), 
         .Z(n7677[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i2_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7646), .D(n7614), 
         .Z(n7677[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i1_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7645), .D(n7613), 
         .Z(n7677[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i15_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7659), .D(n7627), 
         .Z(n7677[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i14_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7658), .D(n7626), 
         .Z(n7677[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i13_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7657), .D(n7625), 
         .Z(n7677[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i12_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7656), .D(n7624), 
         .Z(n7677[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i11_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7655), .D(n7623), 
         .Z(n7677[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3183_i10_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7654), .D(n7622), 
         .Z(n7677[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 n6874_bdd_3_lut_33970 (.A(n7062), .B(\genblk1.ra [9]), .C(n7094), 
         .Z(n40108)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33970.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_33973 (.A(n7140), .B(\genblk1.ra [9]), .C(n7172), 
         .Z(n40109)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33973.init = 16'he2e2;
    LUT4 mux_3183_i9_3_lut_4_lut (.A(n6769), .B(n41382), .C(n7653), .D(n7621), 
         .Z(n7677[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam mux_3183_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 n40169_bdd_3_lut_4_lut (.A(n6766), .B(n41382), .C(n45183), .D(n40169), 
         .Z(n40170)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40169_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n6874_bdd_3_lut_33974 (.A(n7061), .B(\genblk1.ra [9]), .C(n7093), 
         .Z(n40113)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33974.init = 16'he2e2;
    LUT4 n40164_bdd_3_lut_4_lut (.A(n6767), .B(n41382), .C(n45183), .D(n40164), 
         .Z(n40165)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40164_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n6767), .B(n41382), .C(n30012), .D(\write_idx_m[2] ), 
         .Z(n31976)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A !((D)+!C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8070;
    LUT4 i32335_3_lut_4_lut (.A(n6767), .B(n41382), .C(n37504), .D(n37503), 
         .Z(n37507)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32335_3_lut_4_lut.init = 16'hf780;
    LUT4 n6874_bdd_3_lut_33977 (.A(n7139), .B(\genblk1.ra [9]), .C(n7171), 
         .Z(n40114)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33977.init = 16'he2e2;
    LUT4 i32336_3_lut_4_lut (.A(n6767), .B(n41382), .C(n37506), .D(n37505), 
         .Z(n37508)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i32336_3_lut_4_lut.init = 16'hf780;
    LUT4 n6874_bdd_3_lut_33978 (.A(n7060), .B(\genblk1.ra [9]), .C(n7092), 
         .Z(n40118)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33978.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_33981 (.A(n7138), .B(\genblk1.ra [9]), .C(n7170), 
         .Z(n40119)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33981.init = 16'he2e2;
    LUT4 n40227_bdd_3_lut_4_lut (.A(n6751), .B(n41382), .C(n45183), .D(n40227), 
         .Z(n40228)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40227_bdd_3_lut_4_lut.init = 16'h8f80;
    PFUMX i34081 (.BLUT(n40280), .ALUT(n45201), .C0(n45183), .Z(n40281));
    LUT4 n40098_bdd_3_lut_4_lut (.A(n41437), .B(n6781), .C(n45183), .D(n40098), 
         .Z(n40099)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40098_bdd_3_lut_4_lut.init = 16'h2f20;
    LUT4 n6874_bdd_3_lut_33982 (.A(n7059), .B(\genblk1.ra [9]), .C(n7091), 
         .Z(n40123)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33982.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_33985 (.A(n7137), .B(\genblk1.ra [9]), .C(n7169), 
         .Z(n40124)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33985.init = 16'he2e2;
    LUT4 i1_3_lut_4_lut_adj_384 (.A(n6778), .B(n41382), .C(n41364), .D(n41363), 
         .Z(n30820)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_3_lut_4_lut_adj_384.init = 16'hfff8;
    LUT4 n6874_bdd_3_lut_33986 (.A(n7058), .B(\genblk1.ra [9]), .C(n7090), 
         .Z(n40128)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33986.init = 16'he2e2;
    LUT4 i1_2_lut_rep_811_3_lut_4_lut (.A(n6778), .B(n41382), .C(n11834), 
         .D(n41364), .Z(n41216)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_811_3_lut_4_lut.init = 16'hfff8;
    LUT4 n40106_bdd_3_lut_4_lut (.A(n6778), .B(n41382), .C(n45183), .D(n40106), 
         .Z(n40107)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40106_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n6874_bdd_3_lut_33989 (.A(n7136), .B(\genblk1.ra [9]), .C(n7168), 
         .Z(n40129)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33989.init = 16'he2e2;
    LUT4 i1_3_lut_rep_876_4_lut_4_lut (.A(n6778), .B(n41382), .C(n32356), 
         .D(n6780), .Z(n41281)) /* synthesis lut_function=(A (B+(C))+!A (B (C+(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_3_lut_rep_876_4_lut_4_lut.init = 16'hfcf8;
    LUT4 i1_2_lut_rep_824_3_lut_4_lut (.A(n6775), .B(n41382), .C(n41367), 
         .D(n41441), .Z(n41229)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_824_3_lut_4_lut.init = 16'hfff8;
    LUT4 i1_2_lut_rep_822_3_lut_4_lut (.A(n6775), .B(n41382), .C(n41367), 
         .D(n41441), .Z(n41227)) /* synthesis lut_function=(A (B+((D)+!C))+!A ((D)+!C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_822_3_lut_4_lut.init = 16'hff8f;
    LUT4 n6874_bdd_3_lut_33990 (.A(n7057), .B(\genblk1.ra [9]), .C(n7089), 
         .Z(n40133)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33990.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_33993 (.A(n7135), .B(\genblk1.ra [9]), .C(n7167), 
         .Z(n40134)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33993.init = 16'he2e2;
    LUT4 n40121_bdd_3_lut_4_lut (.A(n6775), .B(n41382), .C(n45183), .D(n40121), 
         .Z(n40122)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40121_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i33155_2_lut_3_lut_4_lut_4_lut (.A(n6775), .B(n41382), .C(n41319), 
         .D(n41367), .Z(w_result_sel_mul_d)) /* synthesis lut_function=(!(A (B+!(D))+!A (B (C+!(D))+!B !(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i33155_2_lut_3_lut_4_lut_4_lut.init = 16'h3700;
    LUT4 n6874_bdd_3_lut_33994 (.A(n7056), .B(\genblk1.ra [9]), .C(n7088), 
         .Z(n40138)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33994.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_33997 (.A(n7134), .B(\genblk1.ra [9]), .C(n7166), 
         .Z(n40139)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33997.init = 16'he2e2;
    LUT4 n40116_bdd_3_lut_4_lut (.A(n41381), .B(\genblk1.wait_one_tick_done ), 
         .C(n45183), .D(n40116), .Z(n40117)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40116_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_rep_823_3_lut_4_lut_4_lut (.A(n41381), .B(n45105), .C(n41295), 
         .D(n41451), .Z(n41228)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_823_3_lut_4_lut_4_lut.init = 16'hfff7;
    LUT4 n6874_bdd_3_lut_34001 (.A(n7133), .B(\genblk1.ra [9]), .C(n7165), 
         .Z(n40147)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34001.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_33998 (.A(n7055), .B(\genblk1.ra [9]), .C(n7087), 
         .Z(n40146)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_33998.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_34002 (.A(n7054), .B(\genblk1.ra [9]), .C(n7086), 
         .Z(n40151)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34002.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_34005 (.A(n7132), .B(\genblk1.ra [9]), .C(n7164), 
         .Z(n40152)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34005.init = 16'he2e2;
    PFUMX i34079 (.BLUT(n40278), .ALUT(n40277), .C0(\genblk1.ra [10]), 
          .Z(n40279));
    PFUMX i34076 (.BLUT(n40270), .ALUT(n40268), .C0(n37144), .Z(n40271));
    LUT4 n6874_bdd_3_lut_34006 (.A(n7053), .B(\genblk1.ra [9]), .C(n7085), 
         .Z(n40156)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34006.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_34009 (.A(n7131), .B(\genblk1.ra [9]), .C(n7163), 
         .Z(n40157)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34009.init = 16'he2e2;
    LUT4 n40271_bdd_3_lut_4_lut (.A(n6749), .B(n41382), .C(n45183), .D(n40271), 
         .Z(n40272)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40271_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n40232_bdd_3_lut_4_lut (.A(n6750), .B(n41382), .C(n45183), .D(n40232), 
         .Z(n40233)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40232_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n40222_bdd_3_lut_4_lut (.A(n6752), .B(n41382), .C(n45183), .D(n40222), 
         .Z(n40223)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40222_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n6874_bdd_3_lut_34010 (.A(n7052), .B(\genblk1.ra [9]), .C(n7084), 
         .Z(n40161)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34010.init = 16'he2e2;
    LUT4 n40214_bdd_3_lut_4_lut (.A(n6753), .B(n41382), .C(n45183), .D(n40214), 
         .Z(n40215)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40214_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n40209_bdd_3_lut_4_lut (.A(n6754), .B(n41382), .C(n45183), .D(n40209), 
         .Z(n40210)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40209_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n6874_bdd_3_lut_34013 (.A(n7130), .B(\genblk1.ra [9]), .C(n7162), 
         .Z(n40162)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34013.init = 16'he2e2;
    LUT4 n40204_bdd_3_lut_4_lut (.A(n6755), .B(n41382), .C(n45183), .D(n40204), 
         .Z(n40205)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40204_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n40199_bdd_3_lut_4_lut (.A(n6756), .B(n41382), .C(n45183), .D(n40199), 
         .Z(n40200)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40199_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n40194_bdd_3_lut_4_lut (.A(n6757), .B(n41382), .C(n45183), .D(n40194), 
         .Z(n40195)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40194_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n40189_bdd_3_lut_4_lut (.A(n6758), .B(n41382), .C(n45183), .D(n40189), 
         .Z(n40190)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40189_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n40184_bdd_3_lut_4_lut (.A(n6759), .B(n41382), .C(n45183), .D(n40184), 
         .Z(n40185)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40184_bdd_3_lut_4_lut.init = 16'h8f80;
    PFUMX i34068 (.BLUT(n40237), .ALUT(n45202), .C0(n45183), .Z(n40238));
    LUT4 n6874_bdd_3_lut_34014 (.A(n7051), .B(\genblk1.ra [9]), .C(n7083), 
         .Z(n40166)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34014.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_34017 (.A(n7129), .B(\genblk1.ra [9]), .C(n7161), 
         .Z(n40167)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34017.init = 16'he2e2;
    FD1P3DX pc_d_i2_i3 (.D(pc_f[3]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i3.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i4 (.D(pc_f[4]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i4.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i5 (.D(pc_f[5]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i5.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i6 (.D(pc_f[6]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i6.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i7 (.D(pc_f[7]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i7.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i8 (.D(pc_f[8]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i8.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i9 (.D(pc_f[9]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i9.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i10 (.D(pc_f[10]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i10.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i11 (.D(pc_f[11]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i11.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i12 (.D(pc_f[12]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i12.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i13 (.D(pc_f[13]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i13.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i14 (.D(pc_f[14]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i14.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i15 (.D(pc_f[15]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i15.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i16 (.D(pc_f[16]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i16.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i17 (.D(pc_f[17]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i17.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i18 (.D(pc_f[18]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i18.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i19 (.D(pc_f[19]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i19.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i20 (.D(pc_f[20]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i20.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i21 (.D(pc_f[21]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i21.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i22 (.D(pc_f[22]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i22.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i23 (.D(pc_f[23]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i23.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i24 (.D(pc_f[24]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i24.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i25 (.D(pc_f[25]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i25.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i26 (.D(pc_f[26]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i26.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i27 (.D(pc_f[27]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i27.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i28 (.D(pc_f[28]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i28.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i29 (.D(pc_f[29]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i29.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i30 (.D(pc_f[30]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i30.GSR = "ENABLED";
    FD1P3DX pc_d_i2_i31 (.D(pc_f[31]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_d[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i31.GSR = "ENABLED";
    LUT4 n6874_bdd_3_lut_34018 (.A(n7050), .B(\genblk1.ra [9]), .C(n7082), 
         .Z(n40171)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34018.init = 16'he2e2;
    FD1P3DX pc_x_i2_i3 (.D(pc_d[3]), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i3.GSR = "ENABLED";
    PFUMX i34066 (.BLUT(n40235), .ALUT(n40234), .C0(\genblk1.ra [10]), 
          .Z(n40236));
    FD1S3DX \genblk1.wait_one_tick_done_270_rep_1072  (.D(VCC_net), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n45106)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(418[12] 423[38])
    defparam \genblk1.wait_one_tick_done_270_rep_1072 .GSR = "ENABLED";
    LUT4 n6874_bdd_3_lut_34021 (.A(n7128), .B(\genblk1.ra [9]), .C(n7160), 
         .Z(n40172)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34021.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_34022 (.A(n7049), .B(\genblk1.ra [9]), .C(n7081), 
         .Z(n40176)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34022.init = 16'he2e2;
    FD1S3DX \genblk1.wait_one_tick_done_270_rep_1071  (.D(VCC_net), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(n45105)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=771, LSE_RLINE=790 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(418[12] 423[38])
    defparam \genblk1.wait_one_tick_done_270_rep_1071 .GSR = "ENABLED";
    LUT4 n6874_bdd_3_lut_34025 (.A(n7127), .B(\genblk1.ra [9]), .C(n7159), 
         .Z(n40177)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34025.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_34026 (.A(n7044), .B(\genblk1.ra [9]), .C(n7076), 
         .Z(n40181)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34026.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_34029 (.A(n7122), .B(\genblk1.ra [9]), .C(n7154), 
         .Z(n40182)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34029.init = 16'he2e2;
    FD1P3DX pc_x_i2_i4 (.D(pc_d[4]), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i4.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i5 (.D(pc_d[5]), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i5.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i6 (.D(pc_d[6]), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i6.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i7 (.D(pc_d[7]), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i7.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i8 (.D(pc_d[8]), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i8.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i9 (.D(pc_d[9]), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i9.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i10 (.D(pc_d[10]), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i10.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i11 (.D(pc_d[11]), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i11.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i12 (.D(pc_d[12]), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i12.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i13 (.D(pc_d[13]), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i13.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i14 (.D(pc_d[14]), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i14.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i15 (.D(pc_d[15]), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i15.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i16 (.D(pc_d[16]), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i16.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i17 (.D(pc_d[17]), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i17.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i18 (.D(pc_d[18]), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i18.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i19 (.D(pc_d[19]), .SP(REF_CLK_c_enable_1030), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i19.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i20 (.D(pc_d[20]), .SP(REF_CLK_c_enable_1042), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i20.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i21 (.D(pc_d[21]), .SP(REF_CLK_c_enable_1042), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i21.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i22 (.D(pc_d[22]), .SP(REF_CLK_c_enable_1042), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i22.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i23 (.D(pc_d[23]), .SP(REF_CLK_c_enable_1042), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i23.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i24 (.D(pc_d[24]), .SP(REF_CLK_c_enable_1042), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i24.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i25 (.D(pc_d[25]), .SP(REF_CLK_c_enable_1042), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i25.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i26 (.D(pc_d[26]), .SP(REF_CLK_c_enable_1042), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i26.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i27 (.D(pc_d[27]), .SP(REF_CLK_c_enable_1042), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i27.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i28 (.D(pc_d[28]), .SP(REF_CLK_c_enable_1042), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i28.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i29 (.D(pc_d[29]), .SP(REF_CLK_c_enable_1042), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i29.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i30 (.D(pc_d[30]), .SP(REF_CLK_c_enable_1042), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i30.GSR = "ENABLED";
    FD1P3DX pc_x_i2_i31 (.D(pc_d[31]), .SP(REF_CLK_c_enable_1042), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_x[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i31.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i3 (.D(pc_x[3]), .SP(REF_CLK_c_enable_1050), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i3.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i4 (.D(pc_x[4]), .SP(REF_CLK_c_enable_1050), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i4.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i5 (.D(pc_x[5]), .SP(REF_CLK_c_enable_1050), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i5.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i6 (.D(pc_x[6]), .SP(REF_CLK_c_enable_1050), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i6.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i7 (.D(pc_x[7]), .SP(REF_CLK_c_enable_1050), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i7.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i8 (.D(pc_x[8]), .SP(REF_CLK_c_enable_1050), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i8.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i9 (.D(pc_x[9]), .SP(REF_CLK_c_enable_1050), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i9.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i10 (.D(pc_x[10]), .SP(REF_CLK_c_enable_1050), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i10.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i11 (.D(pc_x[11]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i11.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i12 (.D(pc_x[12]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i12.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i13 (.D(pc_x[13]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i13.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i14 (.D(pc_x[14]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i14.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i15 (.D(pc_x[15]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i15.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i16 (.D(pc_x[16]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i16.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i17 (.D(pc_x[17]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i17.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i18 (.D(pc_x[18]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i18.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i19 (.D(pc_x[19]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i19.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i20 (.D(pc_x[20]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i20.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i21 (.D(pc_x[21]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i21.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i22 (.D(pc_x[22]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i22.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i23 (.D(pc_x[23]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i23.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i24 (.D(pc_x[24]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i24.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i25 (.D(pc_x[25]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i25.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i26 (.D(pc_x[26]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i26.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i27 (.D(pc_x[27]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i27.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i28 (.D(pc_x[28]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i28.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i29 (.D(pc_x[29]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i29.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i30 (.D(pc_x[30]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i30.GSR = "ENABLED";
    FD1P3DX pc_m_i2_i31 (.D(pc_x[31]), .SP(REF_CLK_c_enable_1299), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_m[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i31.GSR = "ENABLED";
    FD1S3DX pc_w_i3 (.D(pc_m[3]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i3.GSR = "ENABLED";
    FD1S3DX pc_w_i4 (.D(pc_m[4]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i4.GSR = "ENABLED";
    FD1S3DX pc_w_i5 (.D(pc_m[5]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i5.GSR = "ENABLED";
    FD1S3DX pc_w_i6 (.D(pc_m[6]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i6.GSR = "ENABLED";
    FD1S3DX pc_w_i7 (.D(pc_m[7]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i7.GSR = "ENABLED";
    FD1S3DX pc_w_i8 (.D(pc_m[8]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i8.GSR = "ENABLED";
    FD1S3DX pc_w_i9 (.D(pc_m[9]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i9.GSR = "ENABLED";
    FD1S3DX pc_w_i10 (.D(pc_m[10]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i10.GSR = "ENABLED";
    FD1S3DX pc_w_i11 (.D(pc_m[11]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i11.GSR = "ENABLED";
    FD1S3DX pc_w_i12 (.D(pc_m[12]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i12.GSR = "ENABLED";
    FD1S3DX pc_w_i13 (.D(pc_m[13]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i13.GSR = "ENABLED";
    FD1S3DX pc_w_i14 (.D(pc_m[14]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i14.GSR = "ENABLED";
    FD1S3DX pc_w_i15 (.D(pc_m[15]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i15.GSR = "ENABLED";
    FD1S3DX pc_w_i16 (.D(pc_m[16]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i16.GSR = "ENABLED";
    FD1S3DX pc_w_i17 (.D(pc_m[17]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i17.GSR = "ENABLED";
    FD1S3DX pc_w_i18 (.D(pc_m[18]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i18.GSR = "ENABLED";
    FD1S3DX pc_w_i19 (.D(pc_m[19]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i19.GSR = "ENABLED";
    FD1S3DX pc_w_i20 (.D(pc_m[20]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i20.GSR = "ENABLED";
    FD1S3DX pc_w_i21 (.D(pc_m[21]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i21.GSR = "ENABLED";
    FD1S3DX pc_w_i22 (.D(pc_m[22]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i22.GSR = "ENABLED";
    FD1S3DX pc_w_i23 (.D(pc_m[23]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i23.GSR = "ENABLED";
    FD1S3DX pc_w_i24 (.D(pc_m[24]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i24.GSR = "ENABLED";
    FD1S3DX pc_w_i25 (.D(pc_m[25]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i25.GSR = "ENABLED";
    FD1S3DX pc_w_i26 (.D(pc_m[26]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i26.GSR = "ENABLED";
    FD1S3DX pc_w_i27 (.D(pc_m[27]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i27.GSR = "ENABLED";
    FD1S3DX pc_w_i28 (.D(pc_m[28]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i28.GSR = "ENABLED";
    FD1S3DX pc_w_i29 (.D(pc_m[29]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i29.GSR = "ENABLED";
    FD1S3DX pc_w_i30 (.D(pc_m[30]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i30.GSR = "ENABLED";
    FD1S3DX pc_w_i31 (.D(pc_m[31]), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(pc_w[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_w_i31.GSR = "ENABLED";
    FD1P3DX restart_address_i3 (.D(restart_address_31__N_1628[1]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i3.GSR = "ENABLED";
    FD1P3DX restart_address_i4 (.D(restart_address_31__N_1628[2]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i4.GSR = "ENABLED";
    FD1P3DX restart_address_i5 (.D(restart_address_31__N_1628[3]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i5.GSR = "ENABLED";
    FD1P3DX restart_address_i6 (.D(restart_address_31__N_1628[4]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i6.GSR = "ENABLED";
    FD1P3DX restart_address_i7 (.D(restart_address_31__N_1628[5]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i7.GSR = "ENABLED";
    FD1P3DX restart_address_i8 (.D(restart_address_31__N_1628[6]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i8.GSR = "ENABLED";
    FD1P3DX restart_address_i9 (.D(restart_address_31__N_1628[7]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i9.GSR = "ENABLED";
    FD1P3DX restart_address_i10 (.D(restart_address_31__N_1628[8]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i10.GSR = "ENABLED";
    FD1P3DX restart_address_i11 (.D(restart_address_31__N_1628[9]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i11.GSR = "ENABLED";
    FD1P3DX restart_address_i12 (.D(restart_address_31__N_1628[10]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i12.GSR = "ENABLED";
    FD1P3DX restart_address_i13 (.D(restart_address_31__N_1628[11]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i13.GSR = "ENABLED";
    FD1P3DX restart_address_i14 (.D(restart_address_31__N_1628[12]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i14.GSR = "ENABLED";
    FD1P3DX restart_address_i15 (.D(restart_address_31__N_1628[13]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i15.GSR = "ENABLED";
    FD1P3DX restart_address_i16 (.D(restart_address_31__N_1628[14]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i16.GSR = "ENABLED";
    FD1P3DX restart_address_i17 (.D(restart_address_31__N_1628[15]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i17.GSR = "ENABLED";
    FD1P3DX restart_address_i18 (.D(restart_address_31__N_1628[16]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i18.GSR = "ENABLED";
    FD1P3DX restart_address_i19 (.D(restart_address_31__N_1628[17]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i19.GSR = "ENABLED";
    FD1P3DX restart_address_i20 (.D(restart_address_31__N_1628[18]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i20.GSR = "ENABLED";
    FD1P3DX restart_address_i21 (.D(restart_address_31__N_1628[19]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i21.GSR = "ENABLED";
    FD1P3DX restart_address_i22 (.D(restart_address_31__N_1628[20]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i22.GSR = "ENABLED";
    FD1P3DX restart_address_i23 (.D(restart_address_31__N_1628[21]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i23.GSR = "ENABLED";
    FD1P3DX restart_address_i24 (.D(restart_address_31__N_1628[22]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i24.GSR = "ENABLED";
    FD1P3DX restart_address_i25 (.D(restart_address_31__N_1628[23]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i25.GSR = "ENABLED";
    FD1P3DX restart_address_i26 (.D(restart_address_31__N_1628[24]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i26.GSR = "ENABLED";
    FD1P3DX restart_address_i27 (.D(restart_address_31__N_1628[25]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i27.GSR = "ENABLED";
    FD1P3DX restart_address_i28 (.D(restart_address_31__N_1628[26]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i28.GSR = "ENABLED";
    FD1P3DX restart_address_i29 (.D(restart_address_31__N_1628[27]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i29.GSR = "ENABLED";
    FD1P3DX restart_address_i30 (.D(restart_address_31__N_1628[28]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i30.GSR = "ENABLED";
    FD1P3DX restart_address_i31 (.D(restart_address_31__N_1628[29]), .SP(REF_CLK_c_enable_1100), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(restart_address[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(625[5] 643[8])
    defparam restart_address_i31.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i1 (.D(SHAREDBUS_DAT_O[1]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i1.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i2 (.D(SHAREDBUS_DAT_O[2]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i2.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i3 (.D(SHAREDBUS_DAT_O[3]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i3.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i4 (.D(SHAREDBUS_DAT_O[4]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i4.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i5 (.D(SHAREDBUS_DAT_O[5]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i5.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i6 (.D(SHAREDBUS_DAT_O[6]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i6.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i7 (.D(SHAREDBUS_DAT_O[7]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i7.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i8 (.D(SHAREDBUS_DAT_O[8]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i8.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i9 (.D(SHAREDBUS_DAT_O[9]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i9.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i10 (.D(SHAREDBUS_DAT_O[10]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i10.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i11 (.D(SHAREDBUS_DAT_O[11]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i11.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i12 (.D(SHAREDBUS_DAT_O[12]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i12.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i13 (.D(SHAREDBUS_DAT_O[13]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i13.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i14 (.D(SHAREDBUS_DAT_O[14]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i14.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i15 (.D(SHAREDBUS_DAT_O[15]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i15.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i16 (.D(SHAREDBUS_DAT_O[16]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i16.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i17 (.D(SHAREDBUS_DAT_O[17]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i17.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i18 (.D(SHAREDBUS_DAT_O[18]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i18.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i19 (.D(SHAREDBUS_DAT_O[19]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i19.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i20 (.D(SHAREDBUS_DAT_O[20]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i20.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i21 (.D(SHAREDBUS_DAT_O[21]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i21.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i22 (.D(SHAREDBUS_DAT_O[22]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i22.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i23 (.D(SHAREDBUS_DAT_O[23]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i23.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i24 (.D(SHAREDBUS_DAT_O[24]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i24.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i25 (.D(SHAREDBUS_DAT_O[25]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i25.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i26 (.D(SHAREDBUS_DAT_O[26]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i26.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i27 (.D(SHAREDBUS_DAT_O[27]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i27.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i28 (.D(SHAREDBUS_DAT_O[28]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i28.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i29 (.D(SHAREDBUS_DAT_O[29]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i29.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i30 (.D(SHAREDBUS_DAT_O[30]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i30.GSR = "ENABLED";
    FD1P3DX icache_refill_data_i0_i31 (.D(SHAREDBUS_DAT_O[31]), .SP(REF_CLK_c_enable_1131), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(icache_refill_data[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam icache_refill_data_i0_i31.GSR = "ENABLED";
    FD1P3DX i_adr_o_i2 (.D(i_adr_o_31__N_1531[2]), .SP(REF_CLK_c_enable_1133), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i2.GSR = "ENABLED";
    PFUMX i34063 (.BLUT(n40231), .ALUT(n40229), .C0(n37144), .Z(n40232));
    LUT4 n6874_bdd_3_lut_34030 (.A(n7043), .B(\genblk1.ra [9]), .C(n7075), 
         .Z(n40186)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34030.init = 16'he2e2;
    PFUMX i34059 (.BLUT(n40226), .ALUT(n40224), .C0(n37144), .Z(n40227));
    FD1P3DX i_adr_o_i3 (.D(i_adr_o_31__N_1531[3]), .SP(REF_CLK_c_enable_1133), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\next_cycle_type[2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i3.GSR = "ENABLED";
    FD1P3DX i_adr_o_i4 (.D(icache_refill_address[4]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i4.GSR = "ENABLED";
    FD1P3DX i_adr_o_i5 (.D(icache_refill_address[5]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[5] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i5.GSR = "ENABLED";
    FD1P3DX i_adr_o_i6 (.D(icache_refill_address[6]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[6] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i6.GSR = "ENABLED";
    FD1P3DX i_adr_o_i7 (.D(icache_refill_address[7]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[7] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i7.GSR = "ENABLED";
    FD1P3DX i_adr_o_i8 (.D(icache_refill_address[8]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[8] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i8.GSR = "ENABLED";
    FD1P3DX i_adr_o_i9 (.D(icache_refill_address[9]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[9] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i9.GSR = "ENABLED";
    FD1P3DX i_adr_o_i10 (.D(icache_refill_address[10]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[10] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i10.GSR = "ENABLED";
    FD1P3DX i_adr_o_i11 (.D(icache_refill_address[11]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[11] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i11.GSR = "ENABLED";
    FD1P3DX i_adr_o_i12 (.D(icache_refill_address[12]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[12] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i12.GSR = "ENABLED";
    FD1P3DX i_adr_o_i13 (.D(icache_refill_address[13]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[13] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i13.GSR = "ENABLED";
    FD1P3DX i_adr_o_i14 (.D(icache_refill_address[14]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[14] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i14.GSR = "ENABLED";
    FD1P3DX i_adr_o_i15 (.D(icache_refill_address[15]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[15] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i15.GSR = "ENABLED";
    FD1P3DX i_adr_o_i16 (.D(icache_refill_address[16]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[16] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i16.GSR = "ENABLED";
    FD1P3DX i_adr_o_i17 (.D(icache_refill_address[17]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[17] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i17.GSR = "ENABLED";
    FD1P3DX i_adr_o_i18 (.D(icache_refill_address[18]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[18] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i18.GSR = "ENABLED";
    FD1P3DX i_adr_o_i19 (.D(icache_refill_address[19]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[19] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i19.GSR = "ENABLED";
    FD1P3DX i_adr_o_i20 (.D(icache_refill_address[20]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[20] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i20.GSR = "ENABLED";
    FD1P3DX i_adr_o_i21 (.D(icache_refill_address[21]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[21] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i21.GSR = "ENABLED";
    FD1P3DX i_adr_o_i22 (.D(icache_refill_address[22]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[22] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i22.GSR = "ENABLED";
    FD1P3DX i_adr_o_i23 (.D(icache_refill_address[23]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[23] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i23.GSR = "ENABLED";
    FD1P3DX i_adr_o_i24 (.D(icache_refill_address[24]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[24] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i24.GSR = "ENABLED";
    FD1P3DX i_adr_o_i25 (.D(icache_refill_address[25]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[25] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i25.GSR = "ENABLED";
    FD1P3DX i_adr_o_i26 (.D(icache_refill_address[26]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[26] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i26.GSR = "ENABLED";
    FD1P3DX i_adr_o_i27 (.D(icache_refill_address[27]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[27] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i27.GSR = "ENABLED";
    FD1P3DX i_adr_o_i28 (.D(icache_refill_address[28]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[28] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i28.GSR = "ENABLED";
    FD1P3DX i_adr_o_i29 (.D(icache_refill_address[29]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[29] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i29.GSR = "ENABLED";
    FD1P3DX i_adr_o_i30 (.D(icache_refill_address[30]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[30] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i30.GSR = "ENABLED";
    FD1P3DX i_adr_o_i31 (.D(icache_refill_address[31]), .SP(REF_CLK_c_enable_1161), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\LM32I_ADR_O[31] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i_adr_o_i31.GSR = "ENABLED";
    FD1P3BX pc_f_i2_i3 (.D(pc_a[3]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(pc_f[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i3.GSR = "ENABLED";
    FD1P3BX pc_f_i2_i4 (.D(pc_a[4]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(pc_f[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i4.GSR = "ENABLED";
    FD1P3BX pc_f_i2_i5 (.D(pc_a[5]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(pc_f[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i5.GSR = "ENABLED";
    FD1P3BX pc_f_i2_i6 (.D(pc_a[6]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(pc_f[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i6.GSR = "ENABLED";
    FD1P3BX pc_f_i2_i7 (.D(pc_a[7]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(pc_f[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i7.GSR = "ENABLED";
    FD1P3BX pc_f_i2_i8 (.D(pc_a[8]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(pc_f[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i8.GSR = "ENABLED";
    FD1P3BX pc_f_i2_i9 (.D(pc_a[9]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(pc_f[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i9.GSR = "ENABLED";
    FD1P3BX pc_f_i2_i10 (.D(pc_a[10]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(pc_f[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i10.GSR = "ENABLED";
    FD1P3BX pc_f_i2_i11 (.D(pc_a[11]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(pc_f[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i11.GSR = "ENABLED";
    FD1P3BX pc_f_i2_i12 (.D(pc_a[12]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(pc_f[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i12.GSR = "ENABLED";
    FD1P3BX pc_f_i2_i13 (.D(pc_a[13]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(pc_f[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i13.GSR = "ENABLED";
    FD1P3BX pc_f_i2_i14 (.D(pc_a[14]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(pc_f[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i14.GSR = "ENABLED";
    FD1P3DX pc_f_i2_i15 (.D(pc_a[15]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_f[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i15.GSR = "ENABLED";
    FD1P3DX pc_f_i2_i16 (.D(pc_a[16]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_f[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i16.GSR = "ENABLED";
    FD1P3DX pc_f_i2_i17 (.D(pc_a[17]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_f[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i17.GSR = "ENABLED";
    FD1P3DX pc_f_i2_i18 (.D(pc_a[18]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_f[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i18.GSR = "ENABLED";
    FD1P3DX pc_f_i2_i19 (.D(pc_a[19]), .SP(REF_CLK_c_enable_1178), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_f[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i19.GSR = "ENABLED";
    FD1P3DX pc_f_i2_i20 (.D(pc_a[20]), .SP(REF_CLK_c_enable_1425), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_f[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i20.GSR = "ENABLED";
    FD1P3DX pc_f_i2_i21 (.D(pc_a[21]), .SP(REF_CLK_c_enable_1425), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_f[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i21.GSR = "ENABLED";
    FD1P3DX pc_f_i2_i22 (.D(pc_a[22]), .SP(REF_CLK_c_enable_1425), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_f[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i22.GSR = "ENABLED";
    FD1P3DX pc_f_i2_i23 (.D(pc_a[23]), .SP(REF_CLK_c_enable_1425), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_f[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i23.GSR = "ENABLED";
    FD1P3DX pc_f_i2_i24 (.D(pc_a[24]), .SP(REF_CLK_c_enable_1425), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_f[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i24.GSR = "ENABLED";
    FD1P3DX pc_f_i2_i25 (.D(pc_a[25]), .SP(REF_CLK_c_enable_1425), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_f[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i25.GSR = "ENABLED";
    FD1P3DX pc_f_i2_i26 (.D(pc_a[26]), .SP(REF_CLK_c_enable_1425), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_f[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i26.GSR = "ENABLED";
    FD1P3DX pc_f_i2_i27 (.D(pc_a[27]), .SP(REF_CLK_c_enable_1425), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_f[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i27.GSR = "ENABLED";
    FD1P3DX pc_f_i2_i28 (.D(pc_a[28]), .SP(REF_CLK_c_enable_1425), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_f[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i28.GSR = "ENABLED";
    FD1P3DX pc_f_i2_i29 (.D(pc_a[29]), .SP(REF_CLK_c_enable_1425), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_f[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i29.GSR = "ENABLED";
    FD1P3DX pc_f_i2_i30 (.D(pc_a[30]), .SP(REF_CLK_c_enable_1425), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_f[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i30.GSR = "ENABLED";
    FD1P3DX pc_f_i2_i31 (.D(pc_a[31]), .SP(REF_CLK_c_enable_1425), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(pc_f[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i31.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_880_3_lut_4_lut_4_lut_4_lut (.A(n45105), .B(n6781), 
         .C(n6777), .D(n6776), .Z(n41285)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_880_3_lut_4_lut_4_lut_4_lut.init = 16'hfdff;
    LUT4 instruction_30__I_0_173_i6_2_lut_rep_843_3_lut_4_lut_4_lut_4_lut (.A(n45105), 
         .B(n6781), .C(n6775), .D(n6776), .Z(n41248)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_30__I_0_173_i6_2_lut_rep_843_3_lut_4_lut_4_lut_4_lut.init = 16'hfdff;
    LUT4 n6874_bdd_3_lut_34033 (.A(n7121), .B(\genblk1.ra [9]), .C(n7153), 
         .Z(n40187)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34033.init = 16'he2e2;
    PFUMX i34055 (.BLUT(n40221), .ALUT(n40219), .C0(n37144), .Z(n40222));
    PFUMX i34051 (.BLUT(n40213), .ALUT(n40211), .C0(n37144), .Z(n40214));
    LUT4 n6874_bdd_3_lut_34034 (.A(n7042), .B(\genblk1.ra [9]), .C(n7074), 
         .Z(n40191)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34034.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_34037 (.A(n7120), .B(\genblk1.ra [9]), .C(n7152), 
         .Z(n40192)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34037.init = 16'he2e2;
    PFUMX i34047 (.BLUT(n40208), .ALUT(n40206), .C0(n37144), .Z(n40209));
    LUT4 n6874_bdd_3_lut_34038 (.A(n7041), .B(\genblk1.ra [9]), .C(n7073), 
         .Z(n40196)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34038.init = 16'he2e2;
    LUT4 i15145_2_lut_rep_976 (.A(n6776), .B(n6781), .Z(n41381)) /* synthesis lut_function=(!((B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i15145_2_lut_rep_976.init = 16'h2222;
    LUT4 i2833_2_lut_rep_962_3_lut (.A(n6776), .B(n6781), .C(n45105), 
         .Z(n41367)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i2833_2_lut_rep_962_3_lut.init = 16'h2020;
    LUT4 i1_4_lut_4_lut_4_lut (.A(n6776), .B(n6781), .C(n32046), .D(n45106), 
         .Z(n30888)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_4_lut_4_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_rep_977 (.A(n45105), .B(n6781), .Z(n41382)) /* synthesis lut_function=(!((B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_977.init = 16'h2222;
    PFUMX i34043 (.BLUT(n40203), .ALUT(n40201), .C0(n37144), .Z(n40204));
    LUT4 i1_2_lut_3_lut_rep_1156 (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n6763), .Z(n45201)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_3_lut_rep_1156.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_rep_1157 (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n6762), .Z(n45202)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_3_lut_rep_1157.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_rep_1159 (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n6761), .Z(n45204)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_3_lut_rep_1159.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_rep_1160 (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n6760), .Z(n45205)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_3_lut_rep_1160.init = 16'h2020;
    LUT4 i1_2_lut_rep_891_3_lut (.A(n45105), .B(n6781), .C(n6780), .Z(n41296)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_891_3_lut.init = 16'h2020;
    LUT4 n6874_bdd_3_lut_34041 (.A(n7119), .B(\genblk1.ra [9]), .C(n7151), 
         .Z(n40197)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34041.init = 16'he2e2;
    LUT4 i1_2_lut_rep_945_3_lut (.A(n45105), .B(n6781), .C(n6770), .Z(n41350)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_945_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_946_3_lut (.A(n45105), .B(n6781), .C(n6772), .Z(n41351)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_946_3_lut.init = 16'h2020;
    PFUMX i34039 (.BLUT(n40198), .ALUT(n40196), .C0(n37144), .Z(n40199));
    LUT4 i1_2_lut_rep_890_3_lut (.A(n45105), .B(n6781), .C(n6777), .Z(n41295)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_890_3_lut.init = 16'h2020;
    LUT4 n6874_bdd_3_lut_34042 (.A(n7040), .B(\genblk1.ra [9]), .C(n7072), 
         .Z(n40201)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34042.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_34045 (.A(n7118), .B(\genblk1.ra [9]), .C(n7150), 
         .Z(n40202)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34045.init = 16'he2e2;
    LUT4 i1_2_lut_rep_842_3_lut_4_lut (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n41419), .D(n6777), .Z(n41247)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_842_3_lut_4_lut.init = 16'h2220;
    LUT4 i1_2_lut_rep_943_3_lut (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n6764), .Z(n41348)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_943_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut (.A(\genblk1.wait_one_tick_done ), .B(n6781), .C(n6760), 
         .Z(\instruction_d[11] )) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_385 (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n6761), .Z(\instruction_d[12] )) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_3_lut_adj_385.init = 16'h2020;
    LUT4 n6874_bdd_3_lut_34046 (.A(n7039), .B(\genblk1.ra [9]), .C(n7071), 
         .Z(n40206)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34046.init = 16'he2e2;
    LUT4 i1_2_lut_3_lut_adj_386 (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n6762), .Z(\instruction_d[13] )) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_3_lut_adj_386.init = 16'h2020;
    LUT4 i1_3_lut_4_lut_else_4_lut_adj_387 (.A(\genblk1.wait_one_tick_done ), 
         .B(n6781), .C(n41208), .D(n6766), .Z(n41465)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_3_lut_4_lut_else_4_lut_adj_387.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_adj_388 (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n6763), .Z(\instruction_d[14] )) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_3_lut_adj_388.init = 16'h2020;
    LUT4 i1_2_lut_rep_947_3_lut (.A(n45105), .B(n6781), .C(n6774), .Z(n41352)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_947_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_948_3_lut (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n6773), .Z(n41353)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_948_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_949_3_lut (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n6771), .Z(n41354)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_949_3_lut.init = 16'h2020;
    LUT4 write_idx_m_4__I_0_793_i2_2_lut_3_lut_4_lut (.A(\genblk1.wait_one_tick_done ), 
         .B(n6781), .C(\write_idx_m[1] ), .D(n6771), .Z(n2_adj_166)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam write_idx_m_4__I_0_793_i2_2_lut_3_lut_4_lut.init = 16'hd2f0;
    LUT4 write_idx_x_4__I_0_791_i2_2_lut_3_lut_4_lut (.A(\genblk1.wait_one_tick_done ), 
         .B(n6781), .C(\write_idx_x[1] ), .D(n6771), .Z(n2_adj_167)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam write_idx_x_4__I_0_791_i2_2_lut_3_lut_4_lut.init = 16'hd2f0;
    LUT4 i1_2_lut_rep_950_3_lut (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n6765), .Z(n41355)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_950_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_951_3_lut (.A(n45105), .B(n6781), .C(n6768), .Z(n41356)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_951_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_952_3_lut (.A(n45105), .B(n6781), .C(n6769), .Z(n41357)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_952_3_lut.init = 16'h2020;
    PFUMX i34035 (.BLUT(n40193), .ALUT(n40191), .C0(n37144), .Z(n40194));
    LUT4 write_idx_m_4__I_0_i5_2_lut_3_lut_4_lut (.A(\genblk1.wait_one_tick_done ), 
         .B(n6781), .C(\write_idx_m[4] ), .D(n6769), .Z(n5)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam write_idx_m_4__I_0_i5_2_lut_3_lut_4_lut.init = 16'hd2f0;
    LUT4 i1_2_lut_rep_953_3_lut (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n6766), .Z(n41358)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_953_3_lut.init = 16'h2020;
    LUT4 write_idx_w_4__I_0_i2_2_lut_3_lut_4_lut (.A(\genblk1.wait_one_tick_done ), 
         .B(n6781), .C(n45099), .D(n6766), .Z(n2_adj_168)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam write_idx_w_4__I_0_i2_2_lut_3_lut_4_lut.init = 16'hd2f0;
    LUT4 n6874_bdd_3_lut_34049 (.A(n7117), .B(\genblk1.ra [9]), .C(n7149), 
         .Z(n40207)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34049.init = 16'he2e2;
    PFUMX i34031 (.BLUT(n40188), .ALUT(n40186), .C0(n37144), .Z(n40189));
    LUT4 write_idx_m_4__I_0_i2_2_lut_rep_877_3_lut_4_lut (.A(\genblk1.wait_one_tick_done ), 
         .B(n6781), .C(\write_idx_m[1] ), .D(n6766), .Z(n41282)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam write_idx_m_4__I_0_i2_2_lut_rep_877_3_lut_4_lut.init = 16'hd2f0;
    LUT4 i1_2_lut_rep_954_3_lut (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n6767), .Z(n41359)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_954_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_956_3_lut (.A(n45105), .B(n6781), .C(n6751), .Z(n41361)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_956_3_lut.init = 16'h2020;
    LUT4 i1_3_lut_rep_958_4_lut (.A(n45105), .B(n6781), .C(n6777), .D(n10475), 
         .Z(n41363)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_3_lut_rep_958_4_lut.init = 16'h2220;
    LUT4 i1_2_lut_rep_960_3_lut (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n6778), .Z(n41365)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_960_3_lut.init = 16'h2020;
    LUT4 n6874_bdd_3_lut_34050 (.A(n7038), .B(\genblk1.ra [9]), .C(n7070), 
         .Z(n40211)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34050.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_34053 (.A(n7116), .B(\genblk1.ra [9]), .C(n7148), 
         .Z(n40212)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34053.init = 16'he2e2;
    LUT4 i1_2_lut_rep_961_3_lut (.A(n45105), .B(n6781), .C(n6775), .Z(n41366)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_961_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_963_3_lut (.A(n45105), .B(n6781), .C(n6749), .Z(n41368)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_963_3_lut.init = 16'h2020;
    PFUMX i34027 (.BLUT(n40183), .ALUT(n40181), .C0(n37144), .Z(n40184));
    LUT4 i1_2_lut_rep_964_3_lut (.A(n45105), .B(n6781), .C(n6750), .Z(n41369)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_964_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_965_3_lut (.A(n45105), .B(n6781), .C(n6752), .Z(n41370)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_965_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_966_3_lut (.A(n45105), .B(n6781), .C(n6753), .Z(n41371)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_966_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_967_3_lut (.A(n45105), .B(n6781), .C(n6754), .Z(n41372)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_967_3_lut.init = 16'h2020;
    LUT4 pc_a_31__I_67_i1_3_lut (.A(pc_a_31__N_1720[0]), .B(restart_address[2]), 
         .C(n41178), .Z(pc_a_31__N_1598[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_968_3_lut (.A(n45105), .B(n6781), .C(n6755), .Z(n41373)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_968_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_969_3_lut (.A(n45105), .B(n6781), .C(n6756), .Z(n41374)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_969_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_970_3_lut (.A(n45105), .B(n6781), .C(n6757), .Z(n41375)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_970_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_971_3_lut (.A(n45105), .B(n6781), .C(n6758), .Z(n41376)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_971_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_972_3_lut (.A(n45105), .B(n6781), .C(n6759), .Z(n41377)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_972_3_lut.init = 16'h2020;
    LUT4 i14767_2_lut_3_lut_4_lut_4_lut (.A(\genblk1.wait_one_tick_done ), 
         .B(n6781), .C(n6775), .D(n6776), .Z(n20031)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i14767_2_lut_3_lut_4_lut_4_lut.init = 16'h2000;
    PFUMX i34023 (.BLUT(n40178), .ALUT(n40176), .C0(n37144), .Z(n40179));
    LUT4 pc_a_31__I_67_i2_3_lut (.A(pc_a_31__N_1720[1]), .B(restart_address[3]), 
         .C(n41178), .Z(pc_a_31__N_1598[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i2_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_67_i4_3_lut (.A(pc_a_31__N_1720[3]), .B(restart_address[5]), 
         .C(n41178), .Z(pc_a_31__N_1598[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i4_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_67_i9_3_lut (.A(pc_a_31__N_1720[8]), .B(restart_address[10]), 
         .C(n41178), .Z(pc_a_31__N_1598[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i9_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_67_i10_3_lut (.A(pc_a_31__N_1720[9]), .B(restart_address[11]), 
         .C(n41178), .Z(pc_a_31__N_1598[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i10_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_67_i11_3_lut (.A(pc_a_31__N_1720[10]), .B(restart_address[12]), 
         .C(n41178), .Z(pc_a_31__N_1598[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i11_3_lut.init = 16'hcaca;
    LUT4 n6874_bdd_3_lut_34057 (.A(n7115), .B(\genblk1.ra [9]), .C(n7147), 
         .Z(n40220)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34057.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_34054 (.A(n7037), .B(\genblk1.ra [9]), .C(n7069), 
         .Z(n40219)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34054.init = 16'he2e2;
    LUT4 pc_a_31__I_67_i12_3_lut (.A(pc_a_31__N_1720[11]), .B(restart_address[13]), 
         .C(n41178), .Z(pc_a_31__N_1598[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i12_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_67_i13_3_lut (.A(pc_a_31__N_1720[12]), .B(restart_address[14]), 
         .C(n41178), .Z(pc_a_31__N_1598[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i13_3_lut.init = 16'hcaca;
    PFUMX i34019 (.BLUT(n40173), .ALUT(n40171), .C0(n37144), .Z(n40174));
    LUT4 pc_a_31__I_67_i14_3_lut (.A(pc_a_31__N_1720[13]), .B(restart_address[15]), 
         .C(n41178), .Z(pc_a_31__N_1598[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i14_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_67_i15_3_lut (.A(pc_a_31__N_1720[14]), .B(restart_address[16]), 
         .C(n41178), .Z(pc_a_31__N_1598[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i15_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_67_i16_3_lut (.A(pc_a_31__N_1720[15]), .B(restart_address[17]), 
         .C(n41178), .Z(pc_a_31__N_1598[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i16_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_67_i17_3_lut (.A(pc_a_31__N_1720[16]), .B(restart_address[18]), 
         .C(n41178), .Z(pc_a_31__N_1598[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i17_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_67_i18_3_lut (.A(pc_a_31__N_1720[17]), .B(restart_address[19]), 
         .C(n41178), .Z(pc_a_31__N_1598[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i18_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_67_i19_3_lut (.A(pc_a_31__N_1720[18]), .B(restart_address[20]), 
         .C(n41178), .Z(pc_a_31__N_1598[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i19_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_67_i20_3_lut (.A(pc_a_31__N_1720[19]), .B(restart_address[21]), 
         .C(n41178), .Z(pc_a_31__N_1598[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i20_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_67_i21_3_lut (.A(pc_a_31__N_1720[20]), .B(restart_address[22]), 
         .C(n41178), .Z(pc_a_31__N_1598[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i21_3_lut.init = 16'hcaca;
    PFUMX i34015 (.BLUT(n40168), .ALUT(n40166), .C0(n37144), .Z(n40169));
    PFUMX i34011 (.BLUT(n40163), .ALUT(n40161), .C0(n37144), .Z(n40164));
    LUT4 n6874_bdd_3_lut_34058 (.A(n7036), .B(\genblk1.ra [9]), .C(n7068), 
         .Z(n40224)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34058.init = 16'he2e2;
    LUT4 pc_a_31__I_67_i22_3_lut (.A(pc_a_31__N_1720[21]), .B(restart_address[23]), 
         .C(n41178), .Z(pc_a_31__N_1598[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i22_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_67_i23_3_lut (.A(pc_a_31__N_1720[22]), .B(restart_address[24]), 
         .C(n41178), .Z(pc_a_31__N_1598[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i23_3_lut.init = 16'hcaca;
    PFUMX i34007 (.BLUT(n40158), .ALUT(n40156), .C0(n37144), .Z(n40159));
    LUT4 n6874_bdd_3_lut_34061 (.A(n7114), .B(\genblk1.ra [9]), .C(n7146), 
         .Z(n40225)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34061.init = 16'he2e2;
    PFUMX i34003 (.BLUT(n40153), .ALUT(n40151), .C0(n37144), .Z(n40154));
    LUT4 pc_a_31__I_67_i24_3_lut (.A(pc_a_31__N_1720[23]), .B(restart_address[25]), 
         .C(n41178), .Z(pc_a_31__N_1598[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i24_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_67_i25_3_lut (.A(pc_a_31__N_1720[24]), .B(restart_address[26]), 
         .C(n41178), .Z(pc_a_31__N_1598[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i25_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_389 (.A(n41179), .B(\extended_immediate[31] ), .C(n2_adj_169), 
         .D(n41291), .Z(n2_adj_170)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(414[8:26])
    defparam i1_4_lut_adj_389.init = 16'ha088;
    LUT4 i1_4_lut_adj_390 (.A(n41179), .B(\extended_immediate[31] ), .C(n2_adj_171), 
         .D(n41291), .Z(n2_adj_172)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(414[8:26])
    defparam i1_4_lut_adj_390.init = 16'ha088;
    LUT4 i1_4_lut_adj_391 (.A(n41179), .B(\extended_immediate[31] ), .C(n2_adj_173), 
         .D(n41291), .Z(n2_adj_174)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(414[8:26])
    defparam i1_4_lut_adj_391.init = 16'ha088;
    LUT4 i1_4_lut_adj_392 (.A(n41179), .B(\extended_immediate[31] ), .C(n2_adj_175), 
         .D(n41291), .Z(n2_adj_176)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(414[8:26])
    defparam i1_4_lut_adj_392.init = 16'ha088;
    PFUMX i33999 (.BLUT(n40148), .ALUT(n40146), .C0(n37144), .Z(n40149));
    LUT4 pc_a_31__I_67_i26_3_lut (.A(pc_a_31__N_1720[25]), .B(restart_address[27]), 
         .C(n41178), .Z(pc_a_31__N_1598[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i26_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_67_i27_3_lut (.A(pc_a_31__N_1720[26]), .B(restart_address[28]), 
         .C(n41178), .Z(pc_a_31__N_1598[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i27_3_lut.init = 16'hcaca;
    PFUMX i33995 (.BLUT(n40140), .ALUT(n40138), .C0(n37144), .Z(n40141));
    LUT4 n6874_bdd_3_lut_34062 (.A(n7035), .B(\genblk1.ra [9]), .C(n7067), 
         .Z(n40229)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34062.init = 16'he2e2;
    LUT4 n6874_bdd_3_lut_34074 (.A(n7113), .B(\genblk1.ra [9]), .C(n7145), 
         .Z(n40230)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34074.init = 16'he2e2;
    PFUMX i33991 (.BLUT(n40135), .ALUT(n40133), .C0(n37144), .Z(n40136));
    LUT4 n7079_bdd_3_lut_34065 (.A(n7157), .B(n7125), .C(\genblk1.ra [9]), 
         .Z(n40234)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n7079_bdd_3_lut_34065.init = 16'hacac;
    LUT4 n7079_bdd_3_lut (.A(n7079), .B(n7047), .C(\genblk1.ra [9]), .Z(n40235)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n7079_bdd_3_lut.init = 16'hacac;
    LUT4 pc_a_31__I_67_i28_3_lut (.A(pc_a_31__N_1720[27]), .B(restart_address[29]), 
         .C(n41178), .Z(pc_a_31__N_1598[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i28_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_67_i29_3_lut (.A(pc_a_31__N_1720[28]), .B(restart_address[30]), 
         .C(n41178), .Z(pc_a_31__N_1598[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i29_3_lut.init = 16'hcaca;
    PFUMX i33987 (.BLUT(n40130), .ALUT(n40128), .C0(n37144), .Z(n40131));
    PFUMX i33983 (.BLUT(n40125), .ALUT(n40123), .C0(n37144), .Z(n40126));
    PFUMX i33979 (.BLUT(n40120), .ALUT(n40118), .C0(n37144), .Z(n40121));
    PFUMX i33975 (.BLUT(n40115), .ALUT(n40113), .C0(n37144), .Z(n40116));
    LUT4 pc_a_31__I_67_i30_3_lut (.A(pc_a_31__N_1720[29]), .B(restart_address[31]), 
         .C(n41178), .Z(pc_a_31__N_1598[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_67_i30_3_lut.init = 16'hcaca;
    PFUMX i33971 (.BLUT(n40110), .ALUT(n40108), .C0(n37144), .Z(n40111));
    LUT4 i1_3_lut_adj_393 (.A(n6772), .B(n6774), .C(n6773), .Z(n31807)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_adj_393.init = 16'hfefe;
    LUT4 i1_4_lut_adj_394 (.A(n41296), .B(n6776), .C(n6775), .D(n6779), 
         .Z(n35314)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C (D)))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_4_lut_adj_394.init = 16'h2080;
    LUT4 i1_4_lut_adj_395 (.A(n41229), .B(n6028), .C(n41232), .D(n35032), 
         .Z(n12412)) /* synthesis lut_function=(A (B)+!A (B ((D)+!C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(730[28:31])
    defparam i1_4_lut_adj_395.init = 16'hcc8c;
    LUT4 n6874_bdd_3_lut (.A(n7112), .B(\genblk1.ra [9]), .C(n7144), .Z(n40269)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut.init = 16'he2e2;
    LUT4 i1_3_lut_4_lut_then_4_lut_adj_396 (.A(\genblk1.wait_one_tick_done ), 
         .B(n6781), .C(n41208), .D(n6762), .Z(n41469)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_3_lut_4_lut_then_4_lut_adj_396.init = 16'h2f0f;
    PFUMX i33967 (.BLUT(n40105), .ALUT(n40103), .C0(n37144), .Z(n40106));
    LUT4 i1_3_lut_4_lut_else_4_lut_adj_397 (.A(\genblk1.wait_one_tick_done ), 
         .B(n6781), .C(n41208), .D(n6767), .Z(n41468)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_3_lut_4_lut_else_4_lut_adj_397.init = 16'h2f0f;
    LUT4 n6874_bdd_3_lut_34075 (.A(n7034), .B(\genblk1.ra [9]), .C(n7066), 
         .Z(n40268)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6874_bdd_3_lut_34075.init = 16'he2e2;
    LUT4 i1_4_lut_adj_398 (.A(dcache_refilling), .B(dcache_refill_request), 
         .C(dcache_restart_request), .D(icache_refill_request), .Z(REF_CLK_c_enable_1100)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;
    defparam i1_4_lut_adj_398.init = 16'hcdcc;
    LUT4 restart_address_31__I_0_i1_3_lut (.A(icache_refill_address[2]), .B(pc_w[2]), 
         .C(dcache_refill_request), .Z(restart_address_31__N_1628[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_399 (.A(n949[0]), .B(n32220), .C(n31750), .D(n30241), 
         .Z(locked_N_493)) /* synthesis lut_function=(A+!((C+!(D))+!B)) */ ;
    defparam i1_4_lut_adj_399.init = 16'haeaa;
    PFUMX i33963 (.BLUT(n40097), .ALUT(n40095), .C0(n37144), .Z(n40098));
    LUT4 i1_4_lut_adj_400 (.A(n35314), .B(n41382), .C(n6778), .D(n6777), 
         .Z(n6028)) /* synthesis lut_function=(!((B (C+(D)))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_4_lut_adj_400.init = 16'h222a;
    PFUMX i33959 (.BLUT(n40092), .ALUT(n40090), .C0(n37144), .Z(n40093));
    LUT4 n7080_bdd_3_lut (.A(n7080), .B(n7048), .C(\genblk1.ra [9]), .Z(n40278)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n7080_bdd_3_lut.init = 16'hacac;
    PFUMX i33956 (.BLUT(n40076), .ALUT(n45204), .C0(n45183), .Z(n40077));
    PFUMX i33954 (.BLUT(n40074), .ALUT(n40073), .C0(\genblk1.ra [10]), 
          .Z(n40075));
    LUT4 n7080_bdd_3_lut_34078 (.A(n7158), .B(n7126), .C(\genblk1.ra [9]), 
         .Z(n40277)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n7080_bdd_3_lut_34078.init = 16'hacac;
    PFUMX i33951 (.BLUT(n40071), .ALUT(n45205), .C0(n45183), .Z(n40072));
    PFUMX i34371 (.BLUT(n41477), .ALUT(n41478), .C0(n6780), .Z(write_idx_d[0]));
    PFUMX i33565 (.BLUT(n38967), .ALUT(n38966), .C0(bus_error_f_N_1884), 
          .Z(REF_CLK_c_enable_129));
    LUT4 i1_3_lut_4_lut_then_4_lut_adj_401 (.A(\genblk1.wait_one_tick_done ), 
         .B(n6781), .C(n41208), .D(n6763), .Z(n41472)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_3_lut_4_lut_then_4_lut_adj_401.init = 16'h2f0f;
    PFUMX i33949 (.BLUT(n40069), .ALUT(n40068), .C0(\genblk1.ra [10]), 
          .Z(n40070));
    LUT4 i1_4_lut_adj_402 (.A(n41380), .B(locked_N_493), .C(LM32D_CYC_O), 
         .D(dcache_refilling), .Z(n30879)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_402.init = 16'h8000;
    LUT4 i1_4_lut_adj_403 (.A(n10485), .B(n41441), .C(n45105), .D(n29933), 
         .Z(n31519)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(460[6:19])
    defparam i1_4_lut_adj_403.init = 16'ha080;
    PFUMX i34369 (.BLUT(n41474), .ALUT(n41475), .C0(n6780), .Z(write_idx_d[4]));
    LUT4 icache_refill_request_I_0_2_lut_rep_1005 (.A(icache_refill_request), 
         .B(icache_refill_ready), .Z(n41410)) /* synthesis lut_function=(!((B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(742[17:84])
    defparam icache_refill_request_I_0_2_lut_rep_1005.init = 16'h2222;
    LUT4 i1_2_lut_rep_911_3_lut (.A(icache_refill_request), .B(icache_refill_ready), 
         .C(bus_error_f_N_1884), .Z(REF_CLK_c_enable_1161)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(742[17:84])
    defparam i1_2_lut_rep_911_3_lut.init = 16'h0202;
    LUT4 i1_2_lut_3_lut_adj_404 (.A(icache_refill_request), .B(icache_refill_ready), 
         .C(bus_error_f_N_1884), .Z(REF_CLK_c_enable_1133)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(742[17:84])
    defparam i1_2_lut_3_lut_adj_404.init = 16'hf2f2;
    LUT4 i1_4_lut_adj_405 (.A(selected[1]), .B(REF_CLK_c_enable_1161), .C(n13990), 
         .D(n32478), .Z(REF_CLK_c_enable_406)) /* synthesis lut_function=(A (B)+!A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_405.init = 16'hdccc;
    LUT4 i1_4_lut_adj_406 (.A(bus_error_f_N_1884), .B(\next_cycle_type[2] ), 
         .C(\LM32I_ADR_O[2] ), .D(selected[0]), .Z(n32478)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_406.init = 16'h8000;
    LUT4 i6993_1_lut (.A(bus_error_f_N_1884), .Z(n9336)) /* synthesis lut_function=(!(A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(698[5] 789[8])
    defparam i6993_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_adj_407 (.A(n6781), .B(n31519), .Z(m_result_sel_shift_d)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(418[12] 423[38])
    defparam i1_2_lut_adj_407.init = 16'hbbbb;
    LUT4 i33324_3_lut_rep_803_4_lut (.A(n41382), .B(n6777), .C(n41381), 
         .D(n30058), .Z(n41208)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i33324_3_lut_rep_803_4_lut.init = 16'h7fff;
    LUT4 n40111_bdd_3_lut_4_lut (.A(n41382), .B(n6777), .C(n45183), .D(n40111), 
         .Z(n40112)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam n40111_bdd_3_lut_4_lut.init = 16'h8f80;
    PFUMX i34367 (.BLUT(n41471), .ALUT(n41472), .C0(n6780), .Z(write_idx_d[3]));
    LUT4 i1_2_lut_rep_1032 (.A(\genblk1.wait_one_tick_done ), .B(n6779), 
         .Z(n41437)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_1032.init = 16'h8888;
    LUT4 i1_2_lut_rep_957_3_lut (.A(\genblk1.wait_one_tick_done ), .B(n6779), 
         .C(n6781), .Z(n41362)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_2_lut_rep_957_3_lut.init = 16'h0808;
    LUT4 i1_4_lut_4_lut_4_lut_adj_408 (.A(\genblk1.wait_one_tick_done ), .B(n6779), 
         .C(n6780), .D(n6781), .Z(n32152)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_4_lut_4_lut_4_lut_adj_408.init = 16'h0020;
    LUT4 i13_4_lut_then_4_lut (.A(selected[1]), .B(selected[0]), .C(LM32D_WE_O), 
         .D(\LM32D_ADR_O[1] ), .Z(n41460)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i13_4_lut_then_4_lut.init = 16'hffdf;
    LUT4 i13_4_lut_else_4_lut (.A(selected[1]), .B(selected[0]), .C(LM32D_WE_O), 
         .D(\LM32D_ADR_O[1] ), .Z(n41459)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i13_4_lut_else_4_lut.init = 16'h2000;
    LUT4 i15148_2_lut_rep_1047 (.A(n6779), .B(n6781), .Z(n41452)) /* synthesis lut_function=(!((B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i15148_2_lut_rep_1047.init = 16'h2222;
    LUT4 i14929_2_lut_rep_836_3_lut_4_lut_4_lut (.A(n6779), .B(n6781), .C(n6778), 
         .D(\genblk1.wait_one_tick_done ), .Z(n41241)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i14929_2_lut_rep_836_3_lut_4_lut_4_lut.init = 16'h2000;
    PFUMX i34365 (.BLUT(n41468), .ALUT(n41469), .C0(n6780), .Z(write_idx_d[2]));
    PFUMX pc_a_31__I_0_i30 (.BLUT(pc_a_31__N_1690[29]), .ALUT(pc_a_31__N_1598[29]), 
          .C0(n37918), .Z(pc_a[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    PFUMX i34363 (.BLUT(n41465), .ALUT(n41466), .C0(n6780), .Z(write_idx_d[1]));
    PFUMX pc_a_31__I_0_i29 (.BLUT(pc_a_31__N_1690[28]), .ALUT(pc_a_31__N_1598[28]), 
          .C0(n37916), .Z(pc_a[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    PFUMX pc_a_31__I_0_i28 (.BLUT(pc_a_31__N_1690[27]), .ALUT(pc_a_31__N_1598[27]), 
          .C0(n37917), .Z(pc_a[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    PFUMX pc_a_31__I_0_i27 (.BLUT(pc_a_31__N_1690[26]), .ALUT(pc_a_31__N_1598[26]), 
          .C0(n37919), .Z(pc_a[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    PFUMX pc_a_31__I_0_i26 (.BLUT(pc_a_31__N_1690[25]), .ALUT(pc_a_31__N_1598[25]), 
          .C0(n37915), .Z(pc_a[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    PFUMX pc_a_31__I_0_i25 (.BLUT(pc_a_31__N_1690[24]), .ALUT(pc_a_31__N_1598[24]), 
          .C0(n37915), .Z(pc_a[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    PFUMX pc_a_31__I_0_i24 (.BLUT(pc_a_31__N_1690[23]), .ALUT(pc_a_31__N_1598[23]), 
          .C0(n37919), .Z(pc_a[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    PFUMX pc_a_31__I_0_i23 (.BLUT(pc_a_31__N_1690[22]), .ALUT(pc_a_31__N_1598[22]), 
          .C0(n37917), .Z(pc_a[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    PFUMX pc_a_31__I_0_i22 (.BLUT(pc_a_31__N_1690[21]), .ALUT(pc_a_31__N_1598[21]), 
          .C0(n37916), .Z(pc_a[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    LUT4 i1_3_lut_4_lut_then_4_lut_adj_409 (.A(\genblk1.wait_one_tick_done ), 
         .B(n6781), .C(n41208), .D(n6761), .Z(n41466)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam i1_3_lut_4_lut_then_4_lut_adj_409.init = 16'h2000;
    LUT4 restart_address_31__I_0_i2_3_lut (.A(icache_refill_address[3]), .B(pc_w[3]), 
         .C(dcache_refill_request), .Z(restart_address_31__N_1628[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 restart_address_31__I_0_i3_3_lut (.A(icache_refill_address[4]), .B(pc_w[4]), 
         .C(dcache_refill_request), .Z(restart_address_31__N_1628[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 restart_address_31__I_0_i4_3_lut (.A(icache_refill_address[5]), .B(pc_w[5]), 
         .C(dcache_refill_request), .Z(restart_address_31__N_1628[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 restart_address_31__I_0_i5_3_lut (.A(icache_refill_address[6]), .B(pc_w[6]), 
         .C(dcache_refill_request), .Z(restart_address_31__N_1628[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i5_3_lut.init = 16'hcaca;
    PFUMX pc_a_31__I_0_i21 (.BLUT(pc_a_31__N_1690[20]), .ALUT(pc_a_31__N_1598[20]), 
          .C0(n37918), .Z(pc_a[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    PFUMX pc_a_31__I_0_i20 (.BLUT(pc_a_31__N_1690[19]), .ALUT(pc_a_31__N_1598[19]), 
          .C0(n37914), .Z(pc_a[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    LUT4 restart_address_31__I_0_i6_3_lut (.A(icache_refill_address[7]), .B(pc_w[7]), 
         .C(dcache_refill_request), .Z(restart_address_31__N_1628[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i6_3_lut.init = 16'hcaca;
    PFUMX pc_a_31__I_0_i19 (.BLUT(pc_a_31__N_1690[18]), .ALUT(pc_a_31__N_1598[18]), 
          .C0(n37914), .Z(pc_a[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    PFUMX pc_a_31__I_0_i18 (.BLUT(pc_a_31__N_1690[17]), .ALUT(pc_a_31__N_1598[17]), 
          .C0(n37915), .Z(pc_a[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    LUT4 restart_address_31__I_0_i7_3_lut (.A(icache_refill_address[8]), .B(pc_w[8]), 
         .C(dcache_refill_request), .Z(restart_address_31__N_1628[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i7_3_lut.init = 16'hcaca;
    PFUMX pc_a_31__I_0_i17 (.BLUT(pc_a_31__N_1690[16]), .ALUT(pc_a_31__N_1598[16]), 
          .C0(n37919), .Z(pc_a[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    LUT4 restart_address_31__I_0_i8_3_lut (.A(icache_refill_address[9]), .B(pc_w[9]), 
         .C(dcache_refill_request), .Z(restart_address_31__N_1628[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i8_3_lut.init = 16'hcaca;
    PFUMX pc_a_31__I_0_i16 (.BLUT(pc_a_31__N_1690[15]), .ALUT(pc_a_31__N_1598[15]), 
          .C0(n37917), .Z(pc_a[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    LUT4 restart_address_31__I_0_i9_3_lut (.A(icache_refill_address[10]), 
         .B(pc_w[10]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i9_3_lut.init = 16'hcaca;
    PFUMX pc_a_31__I_0_i15 (.BLUT(pc_a_31__N_1690[14]), .ALUT(pc_a_31__N_1598[14]), 
          .C0(n37918), .Z(pc_a[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    LUT4 restart_address_31__I_0_i10_3_lut (.A(icache_refill_address[11]), 
         .B(pc_w[11]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i10_3_lut.init = 16'hcaca;
    PFUMX pc_a_31__I_0_i14 (.BLUT(pc_a_31__N_1690[13]), .ALUT(pc_a_31__N_1598[13]), 
          .C0(n36389), .Z(pc_a[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    LUT4 restart_address_31__I_0_i11_3_lut (.A(icache_refill_address[12]), 
         .B(pc_w[12]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 restart_address_31__I_0_i12_3_lut (.A(icache_refill_address[13]), 
         .B(pc_w[13]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i12_3_lut.init = 16'hcaca;
    PFUMX pc_a_31__I_0_i13 (.BLUT(pc_a_31__N_1690[12]), .ALUT(pc_a_31__N_1598[12]), 
          .C0(n37916), .Z(pc_a[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    LUT4 restart_address_31__I_0_i13_3_lut (.A(icache_refill_address[14]), 
         .B(pc_w[14]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i13_3_lut.init = 16'hcaca;
    PFUMX pc_a_31__I_0_i12 (.BLUT(pc_a_31__N_1690[11]), .ALUT(pc_a_31__N_1598[11]), 
          .C0(n37915), .Z(pc_a[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    PFUMX pc_a_31__I_0_i11 (.BLUT(pc_a_31__N_1690[10]), .ALUT(pc_a_31__N_1598[10]), 
          .C0(n37919), .Z(pc_a[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    LUT4 restart_address_31__I_0_i14_3_lut (.A(icache_refill_address[15]), 
         .B(pc_w[15]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i14_3_lut.init = 16'hcaca;
    PFUMX pc_a_31__I_0_i10 (.BLUT(pc_a_31__N_1690[9]), .ALUT(pc_a_31__N_1598[9]), 
          .C0(n37917), .Z(pc_a[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    PFUMX pc_a_31__I_0_i9 (.BLUT(pc_a_31__N_1690[8]), .ALUT(pc_a_31__N_1598[8]), 
          .C0(n37916), .Z(pc_a[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    LUT4 restart_address_31__I_0_i15_3_lut (.A(icache_refill_address[16]), 
         .B(pc_w[16]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i15_3_lut.init = 16'hcaca;
    PFUMX pc_a_31__I_0_i4 (.BLUT(pc_a_31__N_1690[3]), .ALUT(pc_a_31__N_1598[3]), 
          .C0(n37918), .Z(pc_a[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    LUT4 restart_address_31__I_0_i16_3_lut (.A(icache_refill_address[17]), 
         .B(pc_w[17]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i16_3_lut.init = 16'hcaca;
    PFUMX pc_a_31__I_0_i2 (.BLUT(pc_a_31__N_1690[1]), .ALUT(pc_a_31__N_1598[1]), 
          .C0(n37914), .Z(pc_a[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    LUT4 restart_address_31__I_0_i17_3_lut (.A(icache_refill_address[18]), 
         .B(pc_w[18]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i17_3_lut.init = 16'hcaca;
    PFUMX pc_a_31__I_0_i1 (.BLUT(pc_a_31__N_1690[0]), .ALUT(pc_a_31__N_1598[0]), 
          .C0(n37914), .Z(pc_a[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    LUT4 restart_address_31__I_0_i18_3_lut (.A(icache_refill_address[19]), 
         .B(pc_w[19]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i18_3_lut.init = 16'hcaca;
    LUT4 restart_address_31__I_0_i19_3_lut (.A(icache_refill_address[20]), 
         .B(pc_w[20]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i19_3_lut.init = 16'hcaca;
    LUT4 restart_address_31__I_0_i20_3_lut (.A(icache_refill_address[21]), 
         .B(pc_w[21]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i20_3_lut.init = 16'hcaca;
    LUT4 restart_address_31__I_0_i21_3_lut (.A(icache_refill_address[22]), 
         .B(pc_w[22]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i21_3_lut.init = 16'hcaca;
    LUT4 restart_address_31__I_0_i22_3_lut (.A(icache_refill_address[23]), 
         .B(pc_w[23]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i22_3_lut.init = 16'hcaca;
    LUT4 restart_address_31__I_0_i23_3_lut (.A(icache_refill_address[24]), 
         .B(pc_w[24]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i23_3_lut.init = 16'hcaca;
    LUT4 restart_address_31__I_0_i24_3_lut (.A(icache_refill_address[25]), 
         .B(pc_w[25]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i24_3_lut.init = 16'hcaca;
    LUT4 restart_address_31__I_0_i25_3_lut (.A(icache_refill_address[26]), 
         .B(pc_w[26]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i25_3_lut.init = 16'hcaca;
    LUT4 restart_address_31__I_0_i26_3_lut (.A(icache_refill_address[27]), 
         .B(pc_w[27]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i26_3_lut.init = 16'hcaca;
    LUT4 restart_address_31__I_0_i27_3_lut (.A(icache_refill_address[28]), 
         .B(pc_w[28]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i27_3_lut.init = 16'hcaca;
    LUT4 restart_address_31__I_0_i28_3_lut (.A(icache_refill_address[29]), 
         .B(pc_w[29]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i28_3_lut.init = 16'hcaca;
    LUT4 restart_address_31__I_0_i29_3_lut (.A(icache_refill_address[30]), 
         .B(pc_w[30]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i29_3_lut.init = 16'hcaca;
    LUT4 restart_address_31__I_0_i30_3_lut (.A(icache_refill_address[31]), 
         .B(pc_w[31]), .C(dcache_refill_request), .Z(restart_address_31__N_1628[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(631[18] 632[61])
    defparam restart_address_31__I_0_i30_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_410 (.A(bus_error_f_N_1884), .B(n13990), .C(\LM32I_ADR_O[2] ), 
         .D(n41390), .Z(i_adr_o_31__N_1531[2])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_410.init = 16'ha028;
    PFUMX pc_a_31__I_67_i8 (.BLUT(pc_a_31__N_1690[7]), .ALUT(pc_a_31__N_1720[7]), 
          .C0(branch_taken_m), .Z(pc_a_31__N_1598[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    LUT4 i1_4_lut_adj_411 (.A(bus_error_f_N_1884), .B(n1), .C(\next_cycle_type[2] ), 
         .D(n41390), .Z(i_adr_o_31__N_1531[3])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_411.init = 16'ha028;
    LUT4 i1_2_lut_adj_412 (.A(\LM32I_ADR_O[2] ), .B(n13990), .Z(n1)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_412.init = 16'h8888;
    PFUMX pc_a_31__I_67_i7 (.BLUT(pc_a_31__N_1690[6]), .ALUT(pc_a_31__N_1720[6]), 
          .C0(branch_taken_m), .Z(pc_a_31__N_1598[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    PFUMX pc_a_31__I_67_i6 (.BLUT(pc_a_31__N_1690[5]), .ALUT(pc_a_31__N_1720[5]), 
          .C0(branch_taken_m), .Z(pc_a_31__N_1598[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    PFUMX pc_a_31__I_67_i5 (.BLUT(pc_a_31__N_1690[4]), .ALUT(pc_a_31__N_1720[4]), 
          .C0(branch_taken_m), .Z(pc_a_31__N_1598[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    PFUMX pc_a_31__I_67_i3 (.BLUT(pc_a_31__N_1690[2]), .ALUT(pc_a_31__N_1720[2]), 
          .C0(branch_taken_m), .Z(pc_a_31__N_1598[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;
    \lm32_icache(base_address=32'b0,limit=32'b01111111111111111)  icache (.icache_refill_request(icache_refill_request), 
            .REF_CLK_c(REF_CLK_c), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .icache_refill_address({icache_refill_address}), .pc_f({pc_f}), 
            .flush_set({flush_set}), .icache_restart_request(icache_restart_request), 
            .restart_request_N_1998(restart_request_N_1998), .icache_refilling(icache_refilling), 
            .way_match_0__N_2007(way_match_0__N_2007), .\state[2] (\state[2] ), 
            .n41196(n41196), .n15(n15), .q_d(q_d), .n45175(n45175), 
            .valid_x_N_1285(valid_x_N_1285), .n32278(n32278), .n10(n10_adj_177), 
            .n32264(n32264), .n41354(n41354), .n41203(n41203), .n41408(n41408), 
            .n31807(n31807), .flush_set_8__N_1953({flush_set_8__N_1953}), 
            .n9304(n9304), .icache_refill_ready(icache_refill_ready), .n41(n41), 
            .n41187(n41187), .branch_target_d({branch_target_d}), .n157({n157}), 
            .pc_a_31__N_1690({pc_a_31__N_1690}), .n31996(n31996), .cycles_5__N_2934(cycles_5__N_2934), 
            .REF_CLK_c_enable_1366(REF_CLK_c_enable_1366), .REF_CLK_c_enable_1622(REF_CLK_c_enable_1622), 
            .n41172(n41172), .n32618(n32618), .VCC_net(VCC_net), .GND_net(GND_net), 
            .\pc_a[4] (pc_a[4]), .n45183(n45183), .\pc_a[5] (pc_a[5]), 
            .\pc_a[6] (pc_a[6]), .\pc_a[7] (pc_a[7]), .\pc_a[8] (pc_a[8]), 
            .\pc_a[9] (pc_a[9]), .\pc_a[10] (pc_a[10]), .\pc_a[11] (pc_a[11]), 
            .\pc_a[12] (pc_a[12]), .icache_refill_data({icache_refill_data}), 
            .n7066(n7066), .n7067(n7067), .n7068(n7068), .n7069(n7069), 
            .n7070(n7070), .n7071(n7071), .n7072(n7072), .n7073(n7073), 
            .n7074(n7074), .n7075(n7075), .n7076(n7076), .n7077(n7077), 
            .n7078(n7078), .n7079(n7079), .n7080(n7080), .n7081(n7081), 
            .n7082(n7082), .n7083(n7083), .n7084(n7084), .n7085(n7085), 
            .n7086(n7086), .n7087(n7087), .n7088(n7088), .n7089(n7089), 
            .n7090(n7090), .n7091(n7091), .n7092(n7092), .n7093(n7093), 
            .n7094(n7094), .n7095(n7095), .n7096(n7096), .n7097(n7097), 
            .n40162(n40162), .n40163(n40163), .n7144(n7144), .n7145(n7145), 
            .n7146(n7146), .n7147(n7147), .n7148(n7148), .n7149(n7149), 
            .n7150(n7150), .n7151(n7151), .n7152(n7152), .n7153(n7153), 
            .n7154(n7154), .n7155(n7155), .n7156(n7156), .n7157(n7157), 
            .n7158(n7158), .n7159(n7159), .n7160(n7160), .n7161(n7161), 
            .n7162(n7162), .n7163(n7163), .n7164(n7164), .n7165(n7165), 
            .n7166(n7166), .n7167(n7167), .n7168(n7168), .n7169(n7169), 
            .n7170(n7170), .n7171(n7171), .n7172(n7172), .n7173(n7173), 
            .n7174(n7174), .n7175(n7175), .n7112(n7112), .n7113(n7113), 
            .n7114(n7114), .n7115(n7115), .n7116(n7116), .n7117(n7117), 
            .n7118(n7118), .n7119(n7119), .n7120(n7120), .n7121(n7121), 
            .n7122(n7122), .n7123(n7123), .n7124(n7124), .n7125(n7125), 
            .n7126(n7126), .n7127(n7127), .n7128(n7128), .n7129(n7129), 
            .n7130(n7130), .n7131(n7131), .n7132(n7132), .n7133(n7133), 
            .n7134(n7134), .n7135(n7135), .n7136(n7136), .n7137(n7137), 
            .n7138(n7138), .n7139(n7139), .n7140(n7140), .n7141(n7141), 
            .n7142(n7142), .n7143(n7143), .n40157(n40157), .n40158(n40158), 
            .n40152(n40152), .n40153(n40153), .n40147(n40147), .n40148(n40148), 
            .n7034(n7034), .n7035(n7035), .n7036(n7036), .n7037(n7037), 
            .n7038(n7038), .n7039(n7039), .n7040(n7040), .n7041(n7041), 
            .n7042(n7042), .n7043(n7043), .n7044(n7044), .n7045(n7045), 
            .n7046(n7046), .n7047(n7047), .n7048(n7048), .n7049(n7049), 
            .n7050(n7050), .n7051(n7051), .n7052(n7052), .n7053(n7053), 
            .n7054(n7054), .n7055(n7055), .n7056(n7056), .n7057(n7057), 
            .n7058(n7058), .n7059(n7059), .n7060(n7060), .n7061(n7061), 
            .n7062(n7062), .n7063(n7063), .n7064(n7064), .n7065(n7065), 
            .n40139(n40139), .n40140(n40140), .n40134(n40134), .n40135(n40135), 
            .n40129(n40129), .n40130(n40130), .n40124(n40124), .n40125(n40125), 
            .n40119(n40119), .n40120(n40120), .n40114(n40114), .n40115(n40115), 
            .n40109(n40109), .n40110(n40110), .n40104(n40104), .n40105(n40105), 
            .n40096(n40096), .n40097(n40097), .n40091(n40091), .n40092(n40092), 
            .n40269(n40269), .n40270(n40270), .n40070(n40070), .n40071(n40071), 
            .\genblk1.ra[10] (\genblk1.ra [10]), .n37144(n37144), .n40075(n40075), 
            .n40076(n40076), .n40279(n40279), .n40280(n40280), .\pc_a[2] (pc_a[2]), 
            .\pc_a[3] (pc_a[3]), .\genblk1.ra[9] (\genblk1.ra [9]), .REF_CLK_c_enable_1178(REF_CLK_c_enable_1178), 
            .REF_CLK_c_enable_1425(REF_CLK_c_enable_1425), .n40236(n40236), 
            .n40237(n40237), .n40230(n40230), .n40231(n40231), .n40225(n40225), 
            .n40226(n40226), .n40220(n40220), .n40221(n40221), .n40212(n40212), 
            .n40213(n40213), .n40207(n40207), .n40208(n40208), .n40202(n40202), 
            .n40203(n40203), .n40197(n40197), .n40198(n40198), .n40192(n40192), 
            .n40193(n40193), .n40187(n40187), .n40188(n40188), .n40182(n40182), 
            .n40183(n40183), .n40177(n40177), .n40178(n40178), .n40172(n40172), 
            .n40173(n40173), .n40167(n40167), .n40168(n40168)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(443[7] 464[6])
    
endmodule
//
// Verilog Description of module \lm32_icache(base_address=32'b0,limit=32'b01111111111111111) 
//

module \lm32_icache(base_address=32'b0,limit=32'b01111111111111111)  (icache_refill_request, 
            REF_CLK_c, REF_CLK_c_enable_1606, icache_refill_address, pc_f, 
            flush_set, icache_restart_request, restart_request_N_1998, 
            icache_refilling, way_match_0__N_2007, \state[2] , n41196, 
            n15, q_d, n45175, valid_x_N_1285, n32278, n10, n32264, 
            n41354, n41203, n41408, n31807, flush_set_8__N_1953, n9304, 
            icache_refill_ready, n41, n41187, branch_target_d, n157, 
            pc_a_31__N_1690, n31996, cycles_5__N_2934, REF_CLK_c_enable_1366, 
            REF_CLK_c_enable_1622, n41172, n32618, VCC_net, GND_net, 
            \pc_a[4] , n45183, \pc_a[5] , \pc_a[6] , \pc_a[7] , \pc_a[8] , 
            \pc_a[9] , \pc_a[10] , \pc_a[11] , \pc_a[12] , icache_refill_data, 
            n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, 
            n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, 
            n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, 
            n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, 
            n40162, n40163, n7144, n7145, n7146, n7147, n7148, 
            n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, 
            n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, 
            n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, 
            n7173, n7174, n7175, n7112, n7113, n7114, n7115, n7116, 
            n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, 
            n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, 
            n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, 
            n7141, n7142, n7143, n40157, n40158, n40152, n40153, 
            n40147, n40148, n7034, n7035, n7036, n7037, n7038, 
            n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, 
            n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, 
            n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, 
            n7063, n7064, n7065, n40139, n40140, n40134, n40135, 
            n40129, n40130, n40124, n40125, n40119, n40120, n40114, 
            n40115, n40109, n40110, n40104, n40105, n40096, n40097, 
            n40091, n40092, n40269, n40270, n40070, n40071, \genblk1.ra[10] , 
            n37144, n40075, n40076, n40279, n40280, \pc_a[2] , \pc_a[3] , 
            \genblk1.ra[9] , REF_CLK_c_enable_1178, REF_CLK_c_enable_1425, 
            n40236, n40237, n40230, n40231, n40225, n40226, n40220, 
            n40221, n40212, n40213, n40207, n40208, n40202, n40203, 
            n40197, n40198, n40192, n40193, n40187, n40188, n40182, 
            n40183, n40177, n40178, n40172, n40173, n40167, n40168) /* synthesis syn_module_defined=1 */ ;
    output icache_refill_request;
    input REF_CLK_c;
    input REF_CLK_c_enable_1606;
    output [31:2]icache_refill_address;
    input [31:2]pc_f;
    output [8:0]flush_set;
    output icache_restart_request;
    input restart_request_N_1998;
    output icache_refilling;
    output way_match_0__N_2007;
    output \state[2] ;
    input n41196;
    input n15;
    input q_d;
    input n45175;
    output valid_x_N_1285;
    input n32278;
    input n10;
    input n32264;
    input n41354;
    input n41203;
    input n41408;
    input n31807;
    input [8:0]flush_set_8__N_1953;
    output n9304;
    input icache_refill_ready;
    output n41;
    input n41187;
    input [31:2]branch_target_d;
    input [29:0]n157;
    output [29:0]pc_a_31__N_1690;
    input n31996;
    input cycles_5__N_2934;
    output REF_CLK_c_enable_1366;
    output REF_CLK_c_enable_1622;
    input n41172;
    input n32618;
    input VCC_net;
    input GND_net;
    input \pc_a[4] ;
    input n45183;
    input \pc_a[5] ;
    input \pc_a[6] ;
    input \pc_a[7] ;
    input \pc_a[8] ;
    input \pc_a[9] ;
    input \pc_a[10] ;
    input \pc_a[11] ;
    input \pc_a[12] ;
    input [31:0]icache_refill_data;
    output n7066;
    output n7067;
    output n7068;
    output n7069;
    output n7070;
    output n7071;
    output n7072;
    output n7073;
    output n7074;
    output n7075;
    output n7076;
    output n7077;
    output n7078;
    output n7079;
    output n7080;
    output n7081;
    output n7082;
    output n7083;
    output n7084;
    output n7085;
    output n7086;
    output n7087;
    output n7088;
    output n7089;
    output n7090;
    output n7091;
    output n7092;
    output n7093;
    output n7094;
    output n7095;
    output n7096;
    output n7097;
    input n40162;
    output n40163;
    output n7144;
    output n7145;
    output n7146;
    output n7147;
    output n7148;
    output n7149;
    output n7150;
    output n7151;
    output n7152;
    output n7153;
    output n7154;
    output n7155;
    output n7156;
    output n7157;
    output n7158;
    output n7159;
    output n7160;
    output n7161;
    output n7162;
    output n7163;
    output n7164;
    output n7165;
    output n7166;
    output n7167;
    output n7168;
    output n7169;
    output n7170;
    output n7171;
    output n7172;
    output n7173;
    output n7174;
    output n7175;
    output n7112;
    output n7113;
    output n7114;
    output n7115;
    output n7116;
    output n7117;
    output n7118;
    output n7119;
    output n7120;
    output n7121;
    output n7122;
    output n7123;
    output n7124;
    output n7125;
    output n7126;
    output n7127;
    output n7128;
    output n7129;
    output n7130;
    output n7131;
    output n7132;
    output n7133;
    output n7134;
    output n7135;
    output n7136;
    output n7137;
    output n7138;
    output n7139;
    output n7140;
    output n7141;
    output n7142;
    output n7143;
    input n40157;
    output n40158;
    input n40152;
    output n40153;
    input n40147;
    output n40148;
    output n7034;
    output n7035;
    output n7036;
    output n7037;
    output n7038;
    output n7039;
    output n7040;
    output n7041;
    output n7042;
    output n7043;
    output n7044;
    output n7045;
    output n7046;
    output n7047;
    output n7048;
    output n7049;
    output n7050;
    output n7051;
    output n7052;
    output n7053;
    output n7054;
    output n7055;
    output n7056;
    output n7057;
    output n7058;
    output n7059;
    output n7060;
    output n7061;
    output n7062;
    output n7063;
    output n7064;
    output n7065;
    input n40139;
    output n40140;
    input n40134;
    output n40135;
    input n40129;
    output n40130;
    input n40124;
    output n40125;
    input n40119;
    output n40120;
    input n40114;
    output n40115;
    input n40109;
    output n40110;
    input n40104;
    output n40105;
    input n40096;
    output n40097;
    input n40091;
    output n40092;
    input n40269;
    output n40270;
    input n40070;
    output n40071;
    output \genblk1.ra[10] ;
    output n37144;
    input n40075;
    output n40076;
    input n40279;
    output n40280;
    input \pc_a[2] ;
    input \pc_a[3] ;
    output \genblk1.ra[9] ;
    input REF_CLK_c_enable_1178;
    input REF_CLK_c_enable_1425;
    input n40236;
    output n40237;
    input n40230;
    output n40231;
    input n40225;
    output n40226;
    input n40220;
    output n40221;
    input n40212;
    output n40213;
    input n40207;
    output n40208;
    input n40202;
    output n40203;
    input n40197;
    output n40198;
    input n40192;
    output n40193;
    input n40187;
    output n40188;
    input n40182;
    output n40183;
    input n40177;
    output n40178;
    input n40172;
    output n40173;
    input n40167;
    output n40168;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    
    wire n9341, REF_CLK_c_enable_1402;
    wire [8:0]flush_set_8__N_1927;
    wire [10:0]dmem_write_address;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(189[31:49])
    wire [1:0]dmem_write_address_1__N_1919;
    wire [3:0]way_valid;
    
    wire n4, n2, n3, n7490, n7491, n41224, n7486, n7487, n7488, 
        n7489, n30501;
    wire [3:0]state;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(192[26:31])
    
    wire n9345, n9346, n41315, iflush, n32270, n11, n9306, n25, 
        n41171, n7741, n41411;
    wire [3:0]tmem_write_data;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(190[26:41])
    wire [8:0]tmem_write_address;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(187[31:49])
    
    wire way_tag_0__3__N_1918, n35488, n32248, n31939, n35675, n35830, 
        n35681, n32624, n17, n35508, n35506;
    
    FD1S3DX state_FSM_i1 (.D(n9341), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(icache_refill_request));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam state_FSM_i1.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i2 (.D(pc_f[2]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[2])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i2.GSR = "ENABLED";
    FD1S3BX flush_set_i0 (.D(flush_set_8__N_1927[0]), .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), 
            .Q(flush_set[0])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam flush_set_i0.GSR = "ENABLED";
    FD1S3DX refill_offset_i1 (.D(dmem_write_address_1__N_1919[0]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(dmem_write_address[0])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(481[5] 501[8])
    defparam refill_offset_i1.GSR = "ENABLED";
    FD1S3DX restart_request_79 (.D(restart_request_N_1998), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(icache_restart_request)) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam restart_request_79.GSR = "ENABLED";
    FD1S3DX refilling_74 (.D(icache_refill_request), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(icache_refilling)) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(399[9:32])
    defparam refilling_74.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(way_valid[0]), .B(n4), .C(n2), .D(n3), .Z(way_match_0__N_2007)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(303[23:96])
    defparam i1_4_lut.init = 16'hfffd;
    LUT4 way_tag_0__3__I_0_i4_4_lut (.A(n7490), .B(pc_f[15]), .C(n7491), 
         .D(n41224), .Z(n4)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A (B (C (D))+!B !(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(303[23:96])
    defparam way_tag_0__3__I_0_i4_4_lut.init = 16'h3c66;
    LUT4 way_tag_0__3__I_0_i2_4_lut (.A(n7486), .B(pc_f[13]), .C(n7487), 
         .D(n41224), .Z(n2)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A (B (C (D))+!B !(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(303[23:96])
    defparam way_tag_0__3__I_0_i2_4_lut.init = 16'h3c66;
    LUT4 way_tag_0__3__I_0_i3_4_lut (.A(n7488), .B(pc_f[14]), .C(n7489), 
         .D(n41224), .Z(n3)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A (B (C (D))+!B !(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(303[23:96])
    defparam way_tag_0__3__I_0_i3_4_lut.init = 16'h3c66;
    FD1S3DX state_FSM_i2 (.D(n30501), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(\state[2] ));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam state_FSM_i2.GSR = "ENABLED";
    FD1S3DX state_FSM_i3 (.D(n9345), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(state[1]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam state_FSM_i3.GSR = "ENABLED";
    FD1S3BX state_FSM_i4 (.D(n9346), .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), 
            .Q(state[0]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam state_FSM_i4.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i3 (.D(pc_f[3]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[3])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i3.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i4 (.D(pc_f[4]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[4])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i4.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i5 (.D(pc_f[5]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[5])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i5.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i6 (.D(pc_f[6]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[6])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i6.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i7 (.D(pc_f[7]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[7])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i7.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i8 (.D(pc_f[8]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[8])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i8.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i9 (.D(pc_f[9]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[9])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i9.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i10 (.D(pc_f[10]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[10])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i10.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i11 (.D(pc_f[11]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[11])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i11.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i12 (.D(pc_f[12]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[12])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i12.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i13 (.D(pc_f[13]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[13])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i13.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i14 (.D(pc_f[14]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[14])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i14.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i15 (.D(pc_f[15]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[15])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i15.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i16 (.D(pc_f[16]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[16])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i16.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i17 (.D(pc_f[17]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[17])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i17.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i18 (.D(pc_f[18]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[18])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i18.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i19 (.D(pc_f[19]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[19])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i19.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i20 (.D(pc_f[20]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[20])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i20.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i21 (.D(pc_f[21]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[21])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i21.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i22 (.D(pc_f[22]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[22])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i22.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i23 (.D(pc_f[23]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[23])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i23.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i24 (.D(pc_f[24]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[24])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i24.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i25 (.D(pc_f[25]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[25])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i25.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i26 (.D(pc_f[26]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[26])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i26.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i27 (.D(pc_f[27]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[27])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i27.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i28 (.D(pc_f[28]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[28])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i28.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i29 (.D(pc_f[29]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[29])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i29.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i30 (.D(pc_f[30]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[30])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i30.GSR = "ENABLED";
    FD1P3AX refill_address_i2_i31 (.D(pc_f[31]), .SP(REF_CLK_c_enable_1402), 
            .CK(REF_CLK_c), .Q(icache_refill_address[31])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam refill_address_i2_i31.GSR = "ENABLED";
    FD1S3BX flush_set_i1 (.D(flush_set_8__N_1927[1]), .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), 
            .Q(flush_set[1])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam flush_set_i1.GSR = "ENABLED";
    FD1S3BX flush_set_i2 (.D(flush_set_8__N_1927[2]), .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), 
            .Q(flush_set[2])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam flush_set_i2.GSR = "ENABLED";
    FD1S3BX flush_set_i3 (.D(flush_set_8__N_1927[3]), .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), 
            .Q(flush_set[3])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam flush_set_i3.GSR = "ENABLED";
    FD1S3BX flush_set_i4 (.D(flush_set_8__N_1927[4]), .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), 
            .Q(flush_set[4])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam flush_set_i4.GSR = "ENABLED";
    FD1S3BX flush_set_i5 (.D(flush_set_8__N_1927[5]), .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), 
            .Q(flush_set[5])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam flush_set_i5.GSR = "ENABLED";
    FD1S3BX flush_set_i6 (.D(flush_set_8__N_1927[6]), .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), 
            .Q(flush_set[6])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam flush_set_i6.GSR = "ENABLED";
    FD1S3BX flush_set_i7 (.D(flush_set_8__N_1927[7]), .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), 
            .Q(flush_set[7])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam flush_set_i7.GSR = "ENABLED";
    FD1S3BX flush_set_i8 (.D(flush_set_8__N_1927[8]), .CK(REF_CLK_c), .PD(REF_CLK_c_enable_1606), 
            .Q(flush_set[8])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam flush_set_i8.GSR = "ENABLED";
    FD1S3DX refill_offset_i2 (.D(dmem_write_address_1__N_1919[1]), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(dmem_write_address[1])) /* synthesis LSE_LINE_FILE_ID=23, LSE_LCOL=7, LSE_RCOL=6, LSE_LLINE=443, LSE_RLINE=464 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(481[5] 501[8])
    defparam refill_offset_i2.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_363 (.A(n41196), .B(n15), .C(q_d), .D(n45175), 
         .Z(valid_x_N_1285)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_363.init = 16'h1000;
    LUT4 i4051_4_lut (.A(icache_refill_request), .B(n32278), .C(n41315), 
         .D(iflush), .Z(n9341)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A ((D)+!B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam i4051_4_lut.init = 16'h0ace;
    LUT4 i1_2_lut (.A(n32270), .B(n15), .Z(iflush)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut.init = 16'h2222;
    LUT4 i1_4_lut_adj_364 (.A(n41196), .B(n11), .C(n10), .D(n32264), 
         .Z(n32270)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_364.init = 16'h4000;
    LUT4 i1_4_lut_adj_365 (.A(n41354), .B(n41203), .C(n41408), .D(n31807), 
         .Z(n11)) /* synthesis lut_function=(!((B+!(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_365.init = 16'h2022;
    LUT4 select_520_Select_0_i7_4_lut (.A(flush_set[0]), .B(flush_set_8__N_1953[0]), 
         .C(n9306), .D(n9304), .Z(flush_set_8__N_1927[0])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam select_520_Select_0_i7_4_lut.init = 16'heca0;
    LUT4 select_520_Select_0_i5_2_lut (.A(icache_refill_request), .B(\state[2] ), 
         .Z(n9306)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam select_520_Select_0_i5_2_lut.init = 16'heeee;
    LUT4 select_1647_Select_0_i6_2_lut (.A(state[1]), .B(state[0]), .Z(n9304)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam select_1647_Select_0_i6_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_366 (.A(icache_refill_request), .B(dmem_write_address[0]), 
         .C(icache_refill_ready), .D(n25), .Z(dmem_write_address_1__N_1919[0])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A ((D)+!B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(482[9] 500[16])
    defparam i1_4_lut_adj_366.init = 16'h28ec;
    LUT4 i30_3_lut (.A(icache_refill_request), .B(n41171), .C(\state[2] ), 
         .Z(n25)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(482[9] 500[16])
    defparam i30_3_lut.init = 16'hcaca;
    LUT4 select_520_Select_1_i7_4_lut (.A(flush_set[1]), .B(flush_set_8__N_1953[1]), 
         .C(n9306), .D(n9304), .Z(flush_set_8__N_1927[1])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam select_520_Select_1_i7_4_lut.init = 16'heca0;
    LUT4 select_520_Select_2_i7_4_lut (.A(flush_set[2]), .B(flush_set_8__N_1953[2]), 
         .C(n9306), .D(n9304), .Z(flush_set_8__N_1927[2])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam select_520_Select_2_i7_4_lut.init = 16'heca0;
    LUT4 select_520_Select_3_i7_4_lut (.A(flush_set[3]), .B(flush_set_8__N_1953[3]), 
         .C(n9306), .D(n9304), .Z(flush_set_8__N_1927[3])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam select_520_Select_3_i7_4_lut.init = 16'heca0;
    LUT4 select_520_Select_4_i7_4_lut (.A(flush_set[4]), .B(flush_set_8__N_1953[4]), 
         .C(n9306), .D(n9304), .Z(flush_set_8__N_1927[4])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam select_520_Select_4_i7_4_lut.init = 16'heca0;
    LUT4 select_520_Select_5_i7_4_lut (.A(flush_set[5]), .B(flush_set_8__N_1953[5]), 
         .C(n9306), .D(n9304), .Z(flush_set_8__N_1927[5])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam select_520_Select_5_i7_4_lut.init = 16'heca0;
    LUT4 select_520_Select_6_i7_4_lut (.A(flush_set[6]), .B(flush_set_8__N_1953[6]), 
         .C(n9306), .D(n9304), .Z(flush_set_8__N_1927[6])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam select_520_Select_6_i7_4_lut.init = 16'heca0;
    LUT4 select_520_Select_7_i7_4_lut (.A(flush_set[7]), .B(flush_set_8__N_1953[7]), 
         .C(n9306), .D(n9304), .Z(flush_set_8__N_1927[7])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam select_520_Select_7_i7_4_lut.init = 16'heca0;
    LUT4 select_520_Select_8_i7_4_lut (.A(flush_set[8]), .B(flush_set_8__N_1953[8]), 
         .C(n9306), .D(n9304), .Z(flush_set_8__N_1927[8])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam select_520_Select_8_i7_4_lut.init = 16'heca0;
    LUT4 i1_4_lut_adj_367 (.A(icache_refill_request), .B(dmem_write_address[1]), 
         .C(n7741), .D(n25), .Z(dmem_write_address_1__N_1919[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A ((D)+!B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(482[9] 500[16])
    defparam i1_4_lut_adj_367.init = 16'h28ec;
    LUT4 i3279_2_lut (.A(dmem_write_address[0]), .B(icache_refill_ready), 
         .Z(n7741)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(496[13] 497[58])
    defparam i3279_2_lut.init = 16'h8888;
    LUT4 i14787_2_lut_rep_1006 (.A(dmem_write_address[0]), .B(dmem_write_address[1]), 
         .Z(n41411)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14787_2_lut_rep_1006.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut (.A(dmem_write_address[0]), .B(dmem_write_address[1]), 
         .C(icache_restart_request), .D(icache_refill_ready), .Z(n41)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i15454_2_lut_rep_910_3_lut (.A(dmem_write_address[0]), .B(dmem_write_address[1]), 
         .C(icache_refill_ready), .Z(n41315)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15454_2_lut_rep_910_3_lut.init = 16'h8080;
    LUT4 i33104_2_lut_3_lut_4_lut (.A(state[0]), .B(state[1]), .C(dmem_write_address[1]), 
         .D(dmem_write_address[0]), .Z(tmem_write_data[0])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(364[19:30])
    defparam i33104_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 refill_address_12__I_0_i2_3_lut_4_lut (.A(state[0]), .B(state[1]), 
         .C(flush_set[1]), .D(icache_refill_address[5]), .Z(tmem_write_address[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(364[19:30])
    defparam refill_address_12__I_0_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 refill_address_12__I_0_i1_3_lut_4_lut (.A(state[0]), .B(state[1]), 
         .C(flush_set[0]), .D(icache_refill_address[4]), .Z(tmem_write_address[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(364[19:30])
    defparam refill_address_12__I_0_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 refill_address_12__I_0_i7_3_lut_4_lut (.A(state[0]), .B(state[1]), 
         .C(flush_set[6]), .D(icache_refill_address[10]), .Z(tmem_write_address[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(364[19:30])
    defparam refill_address_12__I_0_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 refill_address_12__I_0_i6_3_lut_4_lut (.A(state[0]), .B(state[1]), 
         .C(flush_set[5]), .D(icache_refill_address[9]), .Z(tmem_write_address[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(364[19:30])
    defparam refill_address_12__I_0_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 refill_address_12__I_0_i8_3_lut_4_lut (.A(state[0]), .B(state[1]), 
         .C(flush_set[7]), .D(icache_refill_address[11]), .Z(tmem_write_address[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(364[19:30])
    defparam refill_address_12__I_0_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 refill_address_12__I_0_i9_3_lut_4_lut (.A(state[0]), .B(state[1]), 
         .C(flush_set[8]), .D(icache_refill_address[12]), .Z(tmem_write_address[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(364[19:30])
    defparam refill_address_12__I_0_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 refill_address_12__I_0_i5_3_lut_4_lut (.A(state[0]), .B(state[1]), 
         .C(flush_set[4]), .D(icache_refill_address[8]), .Z(tmem_write_address[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(364[19:30])
    defparam refill_address_12__I_0_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 refill_address_12__I_0_i4_3_lut_4_lut (.A(state[0]), .B(state[1]), 
         .C(flush_set[3]), .D(icache_refill_address[7]), .Z(tmem_write_address[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(364[19:30])
    defparam refill_address_12__I_0_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 refill_address_12__I_0_i3_3_lut_4_lut (.A(state[0]), .B(state[1]), 
         .C(flush_set[2]), .D(icache_refill_address[6]), .Z(tmem_write_address[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(364[19:30])
    defparam refill_address_12__I_0_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 refill_ready_I_0_2_lut_3_lut (.A(state[0]), .B(state[1]), .C(icache_refill_ready), 
         .Z(way_tag_0__3__N_1918)) /* synthesis lut_function=(A+(B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(364[19:30])
    defparam refill_ready_I_0_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut (.A(state[0]), .B(state[1]), .C(flush_set[3]), 
         .Z(n35488)) /* synthesis lut_function=(!(A (C)+!A ((C)+!B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(364[19:30])
    defparam i1_2_lut_3_lut.init = 16'h0e0e;
    LUT4 mux_20_i3_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[4]), .D(n157[2]), .Z(pc_a_31__N_1690[2])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i3_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i5_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[6]), .D(n157[4]), .Z(pc_a_31__N_1690[4])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i5_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i6_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[7]), .D(n157[5]), .Z(pc_a_31__N_1690[5])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i6_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i7_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[8]), .D(n157[6]), .Z(pc_a_31__N_1690[6])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i7_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i8_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[9]), .D(n157[7]), .Z(pc_a_31__N_1690[7])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i8_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i1_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[2]), .D(n157[0]), .Z(pc_a_31__N_1690[0])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i1_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i2_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[3]), .D(n157[1]), .Z(pc_a_31__N_1690[1])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i2_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i4_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[5]), .D(n157[3]), .Z(pc_a_31__N_1690[3])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i4_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i9_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[10]), .D(n157[8]), .Z(pc_a_31__N_1690[8])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i9_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i10_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[11]), .D(n157[9]), .Z(pc_a_31__N_1690[9])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i10_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i11_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[12]), .D(n157[10]), .Z(pc_a_31__N_1690[10])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i11_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i12_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[13]), .D(n157[11]), .Z(pc_a_31__N_1690[11])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i12_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i13_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[14]), .D(n157[12]), .Z(pc_a_31__N_1690[12])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i13_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i14_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[15]), .D(n157[13]), .Z(pc_a_31__N_1690[13])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i14_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i15_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[16]), .D(n157[14]), .Z(pc_a_31__N_1690[14])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i15_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i16_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[17]), .D(n157[15]), .Z(pc_a_31__N_1690[15])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i16_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i17_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[18]), .D(n157[16]), .Z(pc_a_31__N_1690[16])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i17_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i18_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[19]), .D(n157[17]), .Z(pc_a_31__N_1690[17])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i18_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i19_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[20]), .D(n157[18]), .Z(pc_a_31__N_1690[18])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i19_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i20_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[21]), .D(n157[19]), .Z(pc_a_31__N_1690[19])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i20_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i21_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[22]), .D(n157[20]), .Z(pc_a_31__N_1690[20])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i21_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i22_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[23]), .D(n157[21]), .Z(pc_a_31__N_1690[21])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i22_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i23_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[24]), .D(n157[22]), .Z(pc_a_31__N_1690[22])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i23_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i24_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[25]), .D(n157[23]), .Z(pc_a_31__N_1690[23])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i24_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i25_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[26]), .D(n157[24]), .Z(pc_a_31__N_1690[24])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i25_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i26_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[27]), .D(n157[25]), .Z(pc_a_31__N_1690[25])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i26_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i27_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[28]), .D(n157[26]), .Z(pc_a_31__N_1690[26])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i27_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i28_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[29]), .D(n157[27]), .Z(pc_a_31__N_1690[27])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i28_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i29_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[30]), .D(n157[28]), .Z(pc_a_31__N_1690[28])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i29_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_20_i30_4_lut_4_lut (.A(icache_restart_request), .B(n41187), 
         .C(branch_target_d[31]), .D(n157[29]), .Z(pc_a_31__N_1690[29])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(413[5] 469[8])
    defparam mux_20_i30_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i30412_3_lut_rep_766 (.A(n15), .B(n31996), .C(n32270), .Z(n41171)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(448[18] 452[16])
    defparam i30412_3_lut_rep_766.init = 16'h5454;
    LUT4 i994_2_lut_4_lut (.A(n15), .B(n31996), .C(n32270), .D(\state[2] ), 
         .Z(REF_CLK_c_enable_1402)) /* synthesis lut_function=(!(A+!(B (D)+!B (C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(448[18] 452[16])
    defparam i994_2_lut_4_lut.init = 16'h5400;
    LUT4 i951_2_lut_4_lut (.A(n41196), .B(n15), .C(n45175), .D(cycles_5__N_2934), 
         .Z(REF_CLK_c_enable_1366)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i951_2_lut_4_lut.init = 16'h1000;
    LUT4 i2389_2_lut_4_lut (.A(n41196), .B(n15), .C(n45175), .D(n41203), 
         .Z(REF_CLK_c_enable_1622)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;
    defparam i2389_2_lut_4_lut.init = 16'hff10;
    LUT4 i1_4_lut_adj_368 (.A(n32248), .B(iflush), .C(n41172), .D(\state[2] ), 
         .Z(n30501)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam i1_4_lut_adj_368.init = 16'habaa;
    LUT4 i1_4_lut_adj_369 (.A(n31939), .B(icache_refill_request), .C(n41411), 
         .D(icache_refill_ready), .Z(n32248)) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam i1_4_lut_adj_369.init = 16'heaaa;
    LUT4 i1_4_lut_adj_370 (.A(n35675), .B(n35830), .C(n35488), .D(n35681), 
         .Z(n31939)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_370.init = 16'h0010;
    LUT4 i30516_2_lut (.A(flush_set[7]), .B(flush_set[2]), .Z(n35675)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i30516_2_lut.init = 16'heeee;
    LUT4 i30668_4_lut (.A(flush_set[5]), .B(flush_set[1]), .C(flush_set[0]), 
         .D(flush_set[8]), .Z(n35830)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30668_4_lut.init = 16'hfffe;
    LUT4 i30522_2_lut (.A(flush_set[6]), .B(flush_set[4]), .Z(n35681)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i30522_2_lut.init = 16'heeee;
    LUT4 i4055_4_lut (.A(state[1]), .B(n32624), .C(n17), .D(n15), .Z(n9345)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam i4055_4_lut.init = 16'ha0ec;
    LUT4 i1_4_lut_adj_371 (.A(n41196), .B(n11), .C(n10), .D(n32618), 
         .Z(n32624)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_371.init = 16'h4000;
    LUT4 i1_4_lut_adj_372 (.A(n35508), .B(n35506), .C(flush_set[6]), .D(flush_set[2]), 
         .Z(n17)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(419[17:62])
    defparam i1_4_lut_adj_372.init = 16'hfffe;
    LUT4 i1_4_lut_adj_373 (.A(flush_set[3]), .B(flush_set[1]), .C(flush_set[8]), 
         .D(flush_set[4]), .Z(n35508)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(419[17:62])
    defparam i1_4_lut_adj_373.init = 16'hfffe;
    LUT4 i1_3_lut (.A(flush_set[5]), .B(flush_set[0]), .C(flush_set[7]), 
         .Z(n35506)) /* synthesis lut_function=(A+(B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(419[17:62])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i4056_2_lut (.A(state[0]), .B(n17), .Z(n9346)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(414[9] 468[16])
    defparam i4056_2_lut.init = 16'h8888;
    \lm32_ram(data_width=32'sb0100,address_width=32'sb01001)_U3  \memories_0..way_0_tag_ram  (.tmem_write_address({tmem_write_address}), 
            .\tmem_write_data[0] (tmem_write_data[0]), .\icache_refill_address[13] (icache_refill_address[13]), 
            .\icache_refill_address[14] (icache_refill_address[14]), .\icache_refill_address[15] (icache_refill_address[15]), 
            .n7486(n7486), .n7488(n7488), .n7490(n7490), .REF_CLK_c(REF_CLK_c), 
            .way_tag_0__3__N_1918(way_tag_0__3__N_1918), .VCC_net(VCC_net), 
            .GND_net(GND_net), .n7491(n7491), .n7489(n7489), .n7487(n7487), 
            .n41224(n41224), .\way_valid[0] (way_valid[0]), .\pc_a[4] (\pc_a[4] ), 
            .n45183(n45183), .\pc_a[5] (\pc_a[5] ), .\pc_a[6] (\pc_a[6] ), 
            .\pc_a[7] (\pc_a[7] ), .\pc_a[8] (\pc_a[8] ), .\pc_a[9] (\pc_a[9] ), 
            .\pc_a[10] (\pc_a[10] ), .\pc_a[11] (\pc_a[11] ), .\pc_a[12] (\pc_a[12] )) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(276[5] 290[9])
    \lm32_ram(data_width=32,address_width=32'sb01011)  \memories_0..way_0_data_ram  (.REF_CLK_c(REF_CLK_c), 
            .VCC_net(VCC_net), .GND_net(GND_net), .\dmem_write_address[0] (dmem_write_address[0]), 
            .\dmem_write_address[1] (dmem_write_address[1]), .\icache_refill_address[4] (icache_refill_address[4]), 
            .\icache_refill_address[5] (icache_refill_address[5]), .\icache_refill_address[6] (icache_refill_address[6]), 
            .\icache_refill_address[7] (icache_refill_address[7]), .\icache_refill_address[8] (icache_refill_address[8]), 
            .\icache_refill_address[9] (icache_refill_address[9]), .\icache_refill_address[10] (icache_refill_address[10]), 
            .icache_refill_data({icache_refill_data}), .n7066(n7066), .n7067(n7067), 
            .n7068(n7068), .n7069(n7069), .n7070(n7070), .n7071(n7071), 
            .n7072(n7072), .n7073(n7073), .n7074(n7074), .n7075(n7075), 
            .n7076(n7076), .n7077(n7077), .n7078(n7078), .n7079(n7079), 
            .n7080(n7080), .n7081(n7081), .n7082(n7082), .n7083(n7083), 
            .n7084(n7084), .n7085(n7085), .n7086(n7086), .n7087(n7087), 
            .n7088(n7088), .n7089(n7089), .n7090(n7090), .n7091(n7091), 
            .n7092(n7092), .n7093(n7093), .n7094(n7094), .n7095(n7095), 
            .n7096(n7096), .n7097(n7097), .n40162(n40162), .n40163(n40163), 
            .n7144(n7144), .n7145(n7145), .n7146(n7146), .n7147(n7147), 
            .n7148(n7148), .n7149(n7149), .n7150(n7150), .n7151(n7151), 
            .n7152(n7152), .n7153(n7153), .n7154(n7154), .n7155(n7155), 
            .n7156(n7156), .n7157(n7157), .n7158(n7158), .n7159(n7159), 
            .n7160(n7160), .n7161(n7161), .n7162(n7162), .n7163(n7163), 
            .n7164(n7164), .n7165(n7165), .n7166(n7166), .n7167(n7167), 
            .n7168(n7168), .n7169(n7169), .n7170(n7170), .n7171(n7171), 
            .n7172(n7172), .n7173(n7173), .n7174(n7174), .n7175(n7175), 
            .n7112(n7112), .n7113(n7113), .n7114(n7114), .n7115(n7115), 
            .n7116(n7116), .n7117(n7117), .n7118(n7118), .n7119(n7119), 
            .n7120(n7120), .n7121(n7121), .n7122(n7122), .n7123(n7123), 
            .n7124(n7124), .n7125(n7125), .n7126(n7126), .n7127(n7127), 
            .n7128(n7128), .n7129(n7129), .n7130(n7130), .n7131(n7131), 
            .n7132(n7132), .n7133(n7133), .n7134(n7134), .n7135(n7135), 
            .n7136(n7136), .n7137(n7137), .n7138(n7138), .n7139(n7139), 
            .n7140(n7140), .n7141(n7141), .n7142(n7142), .n7143(n7143), 
            .n40157(n40157), .n40158(n40158), .n40152(n40152), .n40153(n40153), 
            .n40147(n40147), .n40148(n40148), .n7034(n7034), .n7035(n7035), 
            .n7036(n7036), .n7037(n7037), .n7038(n7038), .n7039(n7039), 
            .n7040(n7040), .n7041(n7041), .n7042(n7042), .n7043(n7043), 
            .n7044(n7044), .n7045(n7045), .n7046(n7046), .n7047(n7047), 
            .n7048(n7048), .n7049(n7049), .n7050(n7050), .n7051(n7051), 
            .n7052(n7052), .n7053(n7053), .n7054(n7054), .n7055(n7055), 
            .n7056(n7056), .n7057(n7057), .n7058(n7058), .n7059(n7059), 
            .n7060(n7060), .n7061(n7061), .n7062(n7062), .n7063(n7063), 
            .n7064(n7064), .n7065(n7065), .n40139(n40139), .n40140(n40140), 
            .n40134(n40134), .n40135(n40135), .n40129(n40129), .n40130(n40130), 
            .n40124(n40124), .n40125(n40125), .n40119(n40119), .n40120(n40120), 
            .icache_refill_ready(icache_refill_ready), .n40114(n40114), 
            .n40115(n40115), .\icache_refill_address[12] (icache_refill_address[12]), 
            .\icache_refill_address[11] (icache_refill_address[11]), .n40109(n40109), 
            .n40110(n40110), .n40104(n40104), .n40105(n40105), .n40096(n40096), 
            .n40097(n40097), .n40091(n40091), .n40092(n40092), .n40269(n40269), 
            .n40270(n40270), .n40070(n40070), .n40071(n40071), .\genblk1.ra[10] (\genblk1.ra[10] ), 
            .n37144(n37144), .n40075(n40075), .n40076(n40076), .n40279(n40279), 
            .n40280(n40280), .\pc_a[2] (\pc_a[2] ), .n45183(n45183), .\pc_a[3] (\pc_a[3] ), 
            .\pc_a[4] (\pc_a[4] ), .\pc_a[5] (\pc_a[5] ), .\pc_a[6] (\pc_a[6] ), 
            .\pc_a[7] (\pc_a[7] ), .\pc_a[8] (\pc_a[8] ), .\pc_a[9] (\pc_a[9] ), 
            .\pc_a[10] (\pc_a[10] ), .\genblk1.ra[9] (\genblk1.ra[9] ), 
            .REF_CLK_c_enable_1178(REF_CLK_c_enable_1178), .\pc_a[11] (\pc_a[11] ), 
            .REF_CLK_c_enable_1425(REF_CLK_c_enable_1425), .\pc_a[12] (\pc_a[12] ), 
            .n40236(n40236), .n40237(n40237), .n40230(n40230), .n40231(n40231), 
            .n40225(n40225), .n40226(n40226), .n40220(n40220), .n40221(n40221), 
            .n40212(n40212), .n40213(n40213), .n40207(n40207), .n40208(n40208), 
            .n40202(n40202), .n40203(n40203), .n40197(n40197), .n40198(n40198), 
            .n40192(n40192), .n40193(n40193), .n40187(n40187), .n40188(n40188), 
            .n40182(n40182), .n40183(n40183), .n40177(n40177), .n40178(n40178), 
            .n40172(n40172), .n40173(n40173), .n40167(n40167), .n40168(n40168)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_icache.v(239[5] 253[9])
    
endmodule
//
// Verilog Description of module \lm32_ram(data_width=32'sb0100,address_width=32'sb01001)_U3 
//

module \lm32_ram(data_width=32'sb0100,address_width=32'sb01001)_U3  (tmem_write_address, 
            \tmem_write_data[0] , \icache_refill_address[13] , \icache_refill_address[14] , 
            \icache_refill_address[15] , n7486, n7488, n7490, REF_CLK_c, 
            way_tag_0__3__N_1918, VCC_net, GND_net, n7491, n7489, 
            n7487, n41224, \way_valid[0] , \pc_a[4] , n45183, \pc_a[5] , 
            \pc_a[6] , \pc_a[7] , \pc_a[8] , \pc_a[9] , \pc_a[10] , 
            \pc_a[11] , \pc_a[12] ) /* synthesis syn_module_defined=1 */ ;
    input [8:0]tmem_write_address;
    input \tmem_write_data[0] ;
    input \icache_refill_address[13] ;
    input \icache_refill_address[14] ;
    input \icache_refill_address[15] ;
    output n7486;
    output n7488;
    output n7490;
    input REF_CLK_c;
    input way_tag_0__3__N_1918;
    input VCC_net;
    input GND_net;
    output n7491;
    output n7489;
    output n7487;
    output n41224;
    output \way_valid[0] ;
    input \pc_a[4] ;
    input n45183;
    input \pc_a[5] ;
    input \pc_a[6] ;
    input \pc_a[7] ;
    input \pc_a[8] ;
    input \pc_a[9] ;
    input \pc_a[10] ;
    input \pc_a[11] ;
    input \pc_a[12] ;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    wire [8:0]n7452;
    
    wire n7484, n7485, n7482;
    wire [8:0]\genblk1.ra ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(285[31:33])
    
    wire n7479, n7477, n7475, n7473, n7471, n7469, n7467, n7465, 
        n7463, n7481, n27375, n27374;
    
    DP16KD \genblk1.mem0  (.DIA0(\tmem_write_data[0] ), .DIA1(\icache_refill_address[13] ), 
           .DIA2(\icache_refill_address[14] ), .DIA3(\icache_refill_address[15] ), 
           .DIA4(GND_net), .DIA5(GND_net), .DIA6(GND_net), .DIA7(GND_net), 
           .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), .DIA11(GND_net), 
           .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), .DIA15(GND_net), 
           .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), .ADA1(GND_net), 
           .ADA2(tmem_write_address[0]), .ADA3(tmem_write_address[1]), .ADA4(tmem_write_address[2]), 
           .ADA5(tmem_write_address[3]), .ADA6(tmem_write_address[4]), .ADA7(tmem_write_address[5]), 
           .ADA8(tmem_write_address[6]), .ADA9(tmem_write_address[7]), .ADA10(tmem_write_address[8]), 
           .ADA11(GND_net), .ADA12(GND_net), .ADA13(GND_net), .CEA(VCC_net), 
           .OCEA(VCC_net), .CLKA(REF_CLK_c), .WEA(way_tag_0__3__N_1918), 
           .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), 
           .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
           .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
           .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), .DIB11(GND_net), 
           .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), .DIB15(GND_net), 
           .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), .ADB1(GND_net), 
           .ADB2(n7452[0]), .ADB3(n7452[1]), .ADB4(n7452[2]), .ADB5(n7452[3]), 
           .ADB6(n7452[4]), .ADB7(n7452[5]), .ADB8(n7452[6]), .ADB9(n7452[7]), 
           .ADB10(n7452[8]), .ADB11(GND_net), .ADB12(GND_net), .ADB13(GND_net), 
           .CEB(VCC_net), .OCEB(VCC_net), .CLKB(REF_CLK_c), .WEB(GND_net), 
           .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), .RSTB(GND_net), 
           .DOB0(n7484), .DOB1(n7486), .DOB2(n7488), .DOB3(n7490));
    defparam \genblk1.mem0 .DATA_WIDTH_A = 4;
    defparam \genblk1.mem0 .DATA_WIDTH_B = 4;
    defparam \genblk1.mem0 .REGMODE_A = "NOREG";
    defparam \genblk1.mem0 .REGMODE_B = "NOREG";
    defparam \genblk1.mem0 .RESETMODE = "SYNC";
    defparam \genblk1.mem0 .ASYNC_RESET_RELEASE = "SYNC";
    defparam \genblk1.mem0 .WRITEMODE_A = "WRITETHROUGH";
    defparam \genblk1.mem0 .WRITEMODE_B = "WRITETHROUGH";
    defparam \genblk1.mem0 .CSDECODE_A = "0b000";
    defparam \genblk1.mem0 .CSDECODE_B = "0b000";
    defparam \genblk1.mem0 .GSR = "DISABLED";
    defparam \genblk1.mem0 .INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INIT_DATA = "STATIC";
    FD1S3AX \genblk1.mem  (.D(\icache_refill_address[15] ), .CK(REF_CLK_c), 
            .Q(n7491));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3114  (.D(\icache_refill_address[14] ), .CK(REF_CLK_c), 
            .Q(n7489));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3114 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3113  (.D(\icache_refill_address[13] ), .CK(REF_CLK_c), 
            .Q(n7487));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3113 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3112  (.D(\tmem_write_data[0] ), .CK(REF_CLK_c), 
            .Q(n7485));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_3112 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3111  (.D(way_tag_0__3__N_1918), .CK(REF_CLK_c), 
            .Q(n7482));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3111 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3109  (.D(n7452[8]), .CK(REF_CLK_c), .Q(\genblk1.ra [8]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3109 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3107  (.D(tmem_write_address[8]), .CK(REF_CLK_c), 
            .Q(n7479));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3107 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3106  (.D(n7452[7]), .CK(REF_CLK_c), .Q(\genblk1.ra [7]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3106 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3105  (.D(tmem_write_address[7]), .CK(REF_CLK_c), 
            .Q(n7477));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3105 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3104  (.D(n7452[6]), .CK(REF_CLK_c), .Q(\genblk1.ra [6]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3104 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3103  (.D(tmem_write_address[6]), .CK(REF_CLK_c), 
            .Q(n7475));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3103 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3102  (.D(n7452[5]), .CK(REF_CLK_c), .Q(\genblk1.ra [5]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3102 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3101  (.D(tmem_write_address[5]), .CK(REF_CLK_c), 
            .Q(n7473));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3101 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3100  (.D(n7452[4]), .CK(REF_CLK_c), .Q(\genblk1.ra [4]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3100 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3099  (.D(tmem_write_address[4]), .CK(REF_CLK_c), 
            .Q(n7471));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3099 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3098  (.D(n7452[3]), .CK(REF_CLK_c), .Q(\genblk1.ra [3]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3098 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3097  (.D(tmem_write_address[3]), .CK(REF_CLK_c), 
            .Q(n7469));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3097 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3096  (.D(n7452[2]), .CK(REF_CLK_c), .Q(\genblk1.ra [2]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3096 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3095  (.D(tmem_write_address[2]), .CK(REF_CLK_c), 
            .Q(n7467));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3095 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3094  (.D(n7452[1]), .CK(REF_CLK_c), .Q(\genblk1.ra [1]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3094 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3093  (.D(tmem_write_address[1]), .CK(REF_CLK_c), 
            .Q(n7465));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3093 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3092  (.D(n7452[0]), .CK(REF_CLK_c), .Q(\genblk1.ra [0]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_3092 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_3091  (.D(tmem_write_address[0]), .CK(REF_CLK_c), 
            .Q(n7463));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_3091 .GSR = "ENABLED";
    LUT4 i3110_2_lut_rep_819 (.A(n7482), .B(n7481), .Z(n41224)) /* synthesis lut_function=(A (B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam i3110_2_lut_rep_819.init = 16'h8888;
    LUT4 mux_3114_i1_3_lut_4_lut (.A(n7482), .B(n7481), .C(n7485), .D(n7484), 
         .Z(\way_valid[0] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3114_i1_3_lut_4_lut.init = 16'hf780;
    CCU2C equal_3107_9 (.A0(\genblk1.ra [1]), .B0(n7465), .C0(\genblk1.ra [0]), 
          .D0(n7463), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n27375), .S1(n7481));
    defparam equal_3107_9.INIT0 = 16'h9009;
    defparam equal_3107_9.INIT1 = 16'h0000;
    defparam equal_3107_9.INJECT1_0 = "YES";
    defparam equal_3107_9.INJECT1_1 = "NO";
    CCU2C equal_3107_8 (.A0(\genblk1.ra [5]), .B0(n7473), .C0(\genblk1.ra [4]), 
          .D0(n7471), .A1(\genblk1.ra [3]), .B1(n7469), .C1(\genblk1.ra [2]), 
          .D1(n7467), .CIN(n27374), .COUT(n27375));
    defparam equal_3107_8.INIT0 = 16'h9009;
    defparam equal_3107_8.INIT1 = 16'h9009;
    defparam equal_3107_8.INJECT1_0 = "YES";
    defparam equal_3107_8.INJECT1_1 = "YES";
    CCU2C equal_3107_0 (.A0(\genblk1.ra [8]), .B0(n7479), .C0(GND_net), 
          .D0(VCC_net), .A1(\genblk1.ra [7]), .B1(n7477), .C1(\genblk1.ra [6]), 
          .D1(n7475), .COUT(n27374));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam equal_3107_0.INIT0 = 16'h0009;
    defparam equal_3107_0.INIT1 = 16'h9009;
    defparam equal_3107_0.INJECT1_0 = "NO";
    defparam equal_3107_0.INJECT1_1 = "YES";
    LUT4 mux_3089_i1_3_lut (.A(\pc_a[4] ), .B(\genblk1.ra [0]), .C(n45183), 
         .Z(n7452[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3089_i1_3_lut.init = 16'hcaca;
    LUT4 mux_3089_i2_3_lut (.A(\pc_a[5] ), .B(\genblk1.ra [1]), .C(n45183), 
         .Z(n7452[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3089_i2_3_lut.init = 16'hcaca;
    LUT4 mux_3089_i3_3_lut (.A(\pc_a[6] ), .B(\genblk1.ra [2]), .C(n45183), 
         .Z(n7452[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3089_i3_3_lut.init = 16'hcaca;
    LUT4 mux_3089_i4_3_lut (.A(\pc_a[7] ), .B(\genblk1.ra [3]), .C(n45183), 
         .Z(n7452[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3089_i4_3_lut.init = 16'hcaca;
    LUT4 mux_3089_i5_3_lut (.A(\pc_a[8] ), .B(\genblk1.ra [4]), .C(n45183), 
         .Z(n7452[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3089_i5_3_lut.init = 16'hcaca;
    LUT4 mux_3089_i6_3_lut (.A(\pc_a[9] ), .B(\genblk1.ra [5]), .C(n45183), 
         .Z(n7452[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3089_i6_3_lut.init = 16'hcaca;
    LUT4 mux_3089_i7_3_lut (.A(\pc_a[10] ), .B(\genblk1.ra [6]), .C(n45183), 
         .Z(n7452[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3089_i7_3_lut.init = 16'hcaca;
    LUT4 mux_3089_i8_3_lut (.A(\pc_a[11] ), .B(\genblk1.ra [7]), .C(n45183), 
         .Z(n7452[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3089_i8_3_lut.init = 16'hcaca;
    LUT4 mux_3089_i9_3_lut (.A(\pc_a[12] ), .B(\genblk1.ra [8]), .C(n45183), 
         .Z(n7452[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_3089_i9_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module \lm32_ram(data_width=32,address_width=32'sb01011) 
//

module \lm32_ram(data_width=32,address_width=32'sb01011)  (REF_CLK_c, VCC_net, 
            GND_net, \dmem_write_address[0] , \dmem_write_address[1] , 
            \icache_refill_address[4] , \icache_refill_address[5] , \icache_refill_address[6] , 
            \icache_refill_address[7] , \icache_refill_address[8] , \icache_refill_address[9] , 
            \icache_refill_address[10] , icache_refill_data, n7066, n7067, 
            n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, 
            n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, 
            n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, 
            n7092, n7093, n7094, n7095, n7096, n7097, n40162, 
            n40163, n7144, n7145, n7146, n7147, n7148, n7149, 
            n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, 
            n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, 
            n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, 
            n7174, n7175, n7112, n7113, n7114, n7115, n7116, n7117, 
            n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, 
            n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, 
            n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, 
            n7142, n7143, n40157, n40158, n40152, n40153, n40147, 
            n40148, n7034, n7035, n7036, n7037, n7038, n7039, 
            n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, 
            n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, 
            n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, 
            n7064, n7065, n40139, n40140, n40134, n40135, n40129, 
            n40130, n40124, n40125, n40119, n40120, icache_refill_ready, 
            n40114, n40115, \icache_refill_address[12] , \icache_refill_address[11] , 
            n40109, n40110, n40104, n40105, n40096, n40097, n40091, 
            n40092, n40269, n40270, n40070, n40071, \genblk1.ra[10] , 
            n37144, n40075, n40076, n40279, n40280, \pc_a[2] , n45183, 
            \pc_a[3] , \pc_a[4] , \pc_a[5] , \pc_a[6] , \pc_a[7] , 
            \pc_a[8] , \pc_a[9] , \pc_a[10] , \genblk1.ra[9] , REF_CLK_c_enable_1178, 
            \pc_a[11] , REF_CLK_c_enable_1425, \pc_a[12] , n40236, n40237, 
            n40230, n40231, n40225, n40226, n40220, n40221, n40212, 
            n40213, n40207, n40208, n40202, n40203, n40197, n40198, 
            n40192, n40193, n40187, n40188, n40182, n40183, n40177, 
            n40178, n40172, n40173, n40167, n40168) /* synthesis syn_module_defined=1 */ ;
    input REF_CLK_c;
    input VCC_net;
    input GND_net;
    input \dmem_write_address[0] ;
    input \dmem_write_address[1] ;
    input \icache_refill_address[4] ;
    input \icache_refill_address[5] ;
    input \icache_refill_address[6] ;
    input \icache_refill_address[7] ;
    input \icache_refill_address[8] ;
    input \icache_refill_address[9] ;
    input \icache_refill_address[10] ;
    input [31:0]icache_refill_data;
    output n7066;
    output n7067;
    output n7068;
    output n7069;
    output n7070;
    output n7071;
    output n7072;
    output n7073;
    output n7074;
    output n7075;
    output n7076;
    output n7077;
    output n7078;
    output n7079;
    output n7080;
    output n7081;
    output n7082;
    output n7083;
    output n7084;
    output n7085;
    output n7086;
    output n7087;
    output n7088;
    output n7089;
    output n7090;
    output n7091;
    output n7092;
    output n7093;
    output n7094;
    output n7095;
    output n7096;
    output n7097;
    input n40162;
    output n40163;
    output n7144;
    output n7145;
    output n7146;
    output n7147;
    output n7148;
    output n7149;
    output n7150;
    output n7151;
    output n7152;
    output n7153;
    output n7154;
    output n7155;
    output n7156;
    output n7157;
    output n7158;
    output n7159;
    output n7160;
    output n7161;
    output n7162;
    output n7163;
    output n7164;
    output n7165;
    output n7166;
    output n7167;
    output n7168;
    output n7169;
    output n7170;
    output n7171;
    output n7172;
    output n7173;
    output n7174;
    output n7175;
    output n7112;
    output n7113;
    output n7114;
    output n7115;
    output n7116;
    output n7117;
    output n7118;
    output n7119;
    output n7120;
    output n7121;
    output n7122;
    output n7123;
    output n7124;
    output n7125;
    output n7126;
    output n7127;
    output n7128;
    output n7129;
    output n7130;
    output n7131;
    output n7132;
    output n7133;
    output n7134;
    output n7135;
    output n7136;
    output n7137;
    output n7138;
    output n7139;
    output n7140;
    output n7141;
    output n7142;
    output n7143;
    input n40157;
    output n40158;
    input n40152;
    output n40153;
    input n40147;
    output n40148;
    output n7034;
    output n7035;
    output n7036;
    output n7037;
    output n7038;
    output n7039;
    output n7040;
    output n7041;
    output n7042;
    output n7043;
    output n7044;
    output n7045;
    output n7046;
    output n7047;
    output n7048;
    output n7049;
    output n7050;
    output n7051;
    output n7052;
    output n7053;
    output n7054;
    output n7055;
    output n7056;
    output n7057;
    output n7058;
    output n7059;
    output n7060;
    output n7061;
    output n7062;
    output n7063;
    output n7064;
    output n7065;
    input n40139;
    output n40140;
    input n40134;
    output n40135;
    input n40129;
    output n40130;
    input n40124;
    output n40125;
    input n40119;
    output n40120;
    input icache_refill_ready;
    input n40114;
    output n40115;
    input \icache_refill_address[12] ;
    input \icache_refill_address[11] ;
    input n40109;
    output n40110;
    input n40104;
    output n40105;
    input n40096;
    output n40097;
    input n40091;
    output n40092;
    input n40269;
    output n40270;
    input n40070;
    output n40071;
    output \genblk1.ra[10] ;
    output n37144;
    input n40075;
    output n40076;
    input n40279;
    output n40280;
    input \pc_a[2] ;
    input n45183;
    input \pc_a[3] ;
    input \pc_a[4] ;
    input \pc_a[5] ;
    input \pc_a[6] ;
    input \pc_a[7] ;
    input \pc_a[8] ;
    input \pc_a[9] ;
    input \pc_a[10] ;
    output \genblk1.ra[9] ;
    input REF_CLK_c_enable_1178;
    input \pc_a[11] ;
    input REF_CLK_c_enable_1425;
    input \pc_a[12] ;
    input n40236;
    output n40237;
    input n40230;
    output n40231;
    input n40225;
    output n40226;
    input n40220;
    output n40221;
    input n40212;
    output n40213;
    input n40207;
    output n40208;
    input n40202;
    output n40203;
    input n40197;
    output n40198;
    input n40192;
    output n40193;
    input n40187;
    output n40188;
    input n40182;
    output n40183;
    input n40177;
    output n40178;
    input n40172;
    output n40173;
    input n40167;
    output n40168;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    
    wire REF_CLK_c_enable_36;
    wire [10:0]n6837;
    
    wire n6873, n6872, n6912, REF_CLK_c_enable_42, REF_CLK_c_enable_43, 
        n6914, n6916, n6918, REF_CLK_c_enable_44, n6938, n6920, 
        n6936, n6922, n6934, n6932, n6930, n6928, n6926, n6924, 
        n6910, n6908, n6906, n6904, n6902, n6900, n6898, n6896, 
        n6894, n6892, n6890, n6888, n6886, n6884, n6882, n6880, 
        n6878, n6876, n6870, n6868;
    wire [10:0]\genblk1.ra ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(285[31:33])
    
    wire n6866, n6864, n6862, n6860, n6858, n6856, n6854, n6852, 
        n6850, n27352, n27353, n27354;
    
    PDPW16KD \genblk1.mem2  (.DI0(icache_refill_data[0]), .DI1(icache_refill_data[1]), 
            .DI2(icache_refill_data[2]), .DI3(icache_refill_data[3]), .DI4(icache_refill_data[4]), 
            .DI5(icache_refill_data[5]), .DI6(icache_refill_data[6]), .DI7(icache_refill_data[7]), 
            .DI8(icache_refill_data[8]), .DI9(icache_refill_data[9]), .DI10(icache_refill_data[10]), 
            .DI11(icache_refill_data[11]), .DI12(icache_refill_data[12]), 
            .DI13(icache_refill_data[13]), .DI14(icache_refill_data[14]), 
            .DI15(icache_refill_data[15]), .DI16(icache_refill_data[16]), 
            .DI17(icache_refill_data[17]), .DI18(icache_refill_data[18]), 
            .DI19(icache_refill_data[19]), .DI20(icache_refill_data[20]), 
            .DI21(icache_refill_data[21]), .DI22(icache_refill_data[22]), 
            .DI23(icache_refill_data[23]), .DI24(icache_refill_data[24]), 
            .DI25(icache_refill_data[25]), .DI26(icache_refill_data[26]), 
            .DI27(icache_refill_data[27]), .DI28(icache_refill_data[28]), 
            .DI29(icache_refill_data[29]), .DI30(icache_refill_data[30]), 
            .DI31(icache_refill_data[31]), .DI32(GND_net), .DI33(GND_net), 
            .DI34(GND_net), .DI35(GND_net), .ADW0(\dmem_write_address[0] ), 
            .ADW1(\dmem_write_address[1] ), .ADW2(\icache_refill_address[4] ), 
            .ADW3(\icache_refill_address[5] ), .ADW4(\icache_refill_address[6] ), 
            .ADW5(\icache_refill_address[7] ), .ADW6(\icache_refill_address[8] ), 
            .ADW7(\icache_refill_address[9] ), .ADW8(\icache_refill_address[10] ), 
            .BE0(VCC_net), .BE1(VCC_net), .BE2(VCC_net), .BE3(VCC_net), 
            .CEW(REF_CLK_c_enable_36), .CLKW(REF_CLK_c), .CSW0(GND_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(GND_net), .ADR5(n6837[0]), 
            .ADR6(n6837[1]), .ADR7(n6837[2]), .ADR8(n6837[3]), .ADR9(n6837[4]), 
            .ADR10(n6837[5]), .ADR11(n6837[6]), .ADR12(n6837[7]), .ADR13(n6837[8]), 
            .CER(VCC_net), .OCER(VCC_net), .CLKR(REF_CLK_c), .CSR0(GND_net), 
            .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), .DO0(n7084), 
            .DO1(n7085), .DO2(n7086), .DO3(n7087), .DO4(n7088), .DO5(n7089), 
            .DO6(n7090), .DO7(n7091), .DO8(n7092), .DO9(n7093), .DO10(n7094), 
            .DO11(n7095), .DO12(n7096), .DO13(n7097), .DO18(n7066), 
            .DO19(n7067), .DO20(n7068), .DO21(n7069), .DO22(n7070), 
            .DO23(n7071), .DO24(n7072), .DO25(n7073), .DO26(n7074), 
            .DO27(n7075), .DO28(n7076), .DO29(n7077), .DO30(n7078), 
            .DO31(n7079), .DO32(n7080), .DO33(n7081), .DO34(n7082), 
            .DO35(n7083));
    defparam \genblk1.mem2 .DATA_WIDTH_W = 36;
    defparam \genblk1.mem2 .DATA_WIDTH_R = 36;
    defparam \genblk1.mem2 .GSR = "DISABLED";
    defparam \genblk1.mem2 .REGMODE = "NOREG";
    defparam \genblk1.mem2 .RESETMODE = "SYNC";
    defparam \genblk1.mem2 .ASYNC_RESET_RELEASE = "SYNC";
    defparam \genblk1.mem2 .CSDECODE_W = "0b000";
    defparam \genblk1.mem2 .CSDECODE_R = "0b000";
    defparam \genblk1.mem2 .INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem2 .INIT_DATA = "STATIC";
    LUT4 n40162_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6912), .D(n40162), 
         .Z(n40163)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40162_bdd_3_lut_4_lut.init = 16'hf780;
    PDPW16KD \genblk1.mem3  (.DI0(icache_refill_data[0]), .DI1(icache_refill_data[1]), 
            .DI2(icache_refill_data[2]), .DI3(icache_refill_data[3]), .DI4(icache_refill_data[4]), 
            .DI5(icache_refill_data[5]), .DI6(icache_refill_data[6]), .DI7(icache_refill_data[7]), 
            .DI8(icache_refill_data[8]), .DI9(icache_refill_data[9]), .DI10(icache_refill_data[10]), 
            .DI11(icache_refill_data[11]), .DI12(icache_refill_data[12]), 
            .DI13(icache_refill_data[13]), .DI14(icache_refill_data[14]), 
            .DI15(icache_refill_data[15]), .DI16(icache_refill_data[16]), 
            .DI17(icache_refill_data[17]), .DI18(icache_refill_data[18]), 
            .DI19(icache_refill_data[19]), .DI20(icache_refill_data[20]), 
            .DI21(icache_refill_data[21]), .DI22(icache_refill_data[22]), 
            .DI23(icache_refill_data[23]), .DI24(icache_refill_data[24]), 
            .DI25(icache_refill_data[25]), .DI26(icache_refill_data[26]), 
            .DI27(icache_refill_data[27]), .DI28(icache_refill_data[28]), 
            .DI29(icache_refill_data[29]), .DI30(icache_refill_data[30]), 
            .DI31(icache_refill_data[31]), .DI32(GND_net), .DI33(GND_net), 
            .DI34(GND_net), .DI35(GND_net), .ADW0(\dmem_write_address[0] ), 
            .ADW1(\dmem_write_address[1] ), .ADW2(\icache_refill_address[4] ), 
            .ADW3(\icache_refill_address[5] ), .ADW4(\icache_refill_address[6] ), 
            .ADW5(\icache_refill_address[7] ), .ADW6(\icache_refill_address[8] ), 
            .ADW7(\icache_refill_address[9] ), .ADW8(\icache_refill_address[10] ), 
            .BE0(VCC_net), .BE1(VCC_net), .BE2(VCC_net), .BE3(VCC_net), 
            .CEW(REF_CLK_c_enable_42), .CLKW(REF_CLK_c), .CSW0(GND_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(GND_net), .ADR5(n6837[0]), 
            .ADR6(n6837[1]), .ADR7(n6837[2]), .ADR8(n6837[3]), .ADR9(n6837[4]), 
            .ADR10(n6837[5]), .ADR11(n6837[6]), .ADR12(n6837[7]), .ADR13(n6837[8]), 
            .CER(VCC_net), .OCER(VCC_net), .CLKR(REF_CLK_c), .CSR0(GND_net), 
            .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), .DO0(n7162), 
            .DO1(n7163), .DO2(n7164), .DO3(n7165), .DO4(n7166), .DO5(n7167), 
            .DO6(n7168), .DO7(n7169), .DO8(n7170), .DO9(n7171), .DO10(n7172), 
            .DO11(n7173), .DO12(n7174), .DO13(n7175), .DO18(n7144), 
            .DO19(n7145), .DO20(n7146), .DO21(n7147), .DO22(n7148), 
            .DO23(n7149), .DO24(n7150), .DO25(n7151), .DO26(n7152), 
            .DO27(n7153), .DO28(n7154), .DO29(n7155), .DO30(n7156), 
            .DO31(n7157), .DO32(n7158), .DO33(n7159), .DO34(n7160), 
            .DO35(n7161));
    defparam \genblk1.mem3 .DATA_WIDTH_W = 36;
    defparam \genblk1.mem3 .DATA_WIDTH_R = 36;
    defparam \genblk1.mem3 .GSR = "DISABLED";
    defparam \genblk1.mem3 .REGMODE = "NOREG";
    defparam \genblk1.mem3 .RESETMODE = "SYNC";
    defparam \genblk1.mem3 .ASYNC_RESET_RELEASE = "SYNC";
    defparam \genblk1.mem3 .CSDECODE_W = "0b000";
    defparam \genblk1.mem3 .CSDECODE_R = "0b000";
    defparam \genblk1.mem3 .INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem3 .INIT_DATA = "STATIC";
    PDPW16KD \genblk1.mem1  (.DI0(icache_refill_data[0]), .DI1(icache_refill_data[1]), 
            .DI2(icache_refill_data[2]), .DI3(icache_refill_data[3]), .DI4(icache_refill_data[4]), 
            .DI5(icache_refill_data[5]), .DI6(icache_refill_data[6]), .DI7(icache_refill_data[7]), 
            .DI8(icache_refill_data[8]), .DI9(icache_refill_data[9]), .DI10(icache_refill_data[10]), 
            .DI11(icache_refill_data[11]), .DI12(icache_refill_data[12]), 
            .DI13(icache_refill_data[13]), .DI14(icache_refill_data[14]), 
            .DI15(icache_refill_data[15]), .DI16(icache_refill_data[16]), 
            .DI17(icache_refill_data[17]), .DI18(icache_refill_data[18]), 
            .DI19(icache_refill_data[19]), .DI20(icache_refill_data[20]), 
            .DI21(icache_refill_data[21]), .DI22(icache_refill_data[22]), 
            .DI23(icache_refill_data[23]), .DI24(icache_refill_data[24]), 
            .DI25(icache_refill_data[25]), .DI26(icache_refill_data[26]), 
            .DI27(icache_refill_data[27]), .DI28(icache_refill_data[28]), 
            .DI29(icache_refill_data[29]), .DI30(icache_refill_data[30]), 
            .DI31(icache_refill_data[31]), .DI32(GND_net), .DI33(GND_net), 
            .DI34(GND_net), .DI35(GND_net), .ADW0(\dmem_write_address[0] ), 
            .ADW1(\dmem_write_address[1] ), .ADW2(\icache_refill_address[4] ), 
            .ADW3(\icache_refill_address[5] ), .ADW4(\icache_refill_address[6] ), 
            .ADW5(\icache_refill_address[7] ), .ADW6(\icache_refill_address[8] ), 
            .ADW7(\icache_refill_address[9] ), .ADW8(\icache_refill_address[10] ), 
            .BE0(VCC_net), .BE1(VCC_net), .BE2(VCC_net), .BE3(VCC_net), 
            .CEW(REF_CLK_c_enable_43), .CLKW(REF_CLK_c), .CSW0(GND_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(GND_net), .ADR5(n6837[0]), 
            .ADR6(n6837[1]), .ADR7(n6837[2]), .ADR8(n6837[3]), .ADR9(n6837[4]), 
            .ADR10(n6837[5]), .ADR11(n6837[6]), .ADR12(n6837[7]), .ADR13(n6837[8]), 
            .CER(VCC_net), .OCER(VCC_net), .CLKR(REF_CLK_c), .CSR0(GND_net), 
            .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), .DO0(n7130), 
            .DO1(n7131), .DO2(n7132), .DO3(n7133), .DO4(n7134), .DO5(n7135), 
            .DO6(n7136), .DO7(n7137), .DO8(n7138), .DO9(n7139), .DO10(n7140), 
            .DO11(n7141), .DO12(n7142), .DO13(n7143), .DO18(n7112), 
            .DO19(n7113), .DO20(n7114), .DO21(n7115), .DO22(n7116), 
            .DO23(n7117), .DO24(n7118), .DO25(n7119), .DO26(n7120), 
            .DO27(n7121), .DO28(n7122), .DO29(n7123), .DO30(n7124), 
            .DO31(n7125), .DO32(n7126), .DO33(n7127), .DO34(n7128), 
            .DO35(n7129));
    defparam \genblk1.mem1 .DATA_WIDTH_W = 36;
    defparam \genblk1.mem1 .DATA_WIDTH_R = 36;
    defparam \genblk1.mem1 .GSR = "DISABLED";
    defparam \genblk1.mem1 .REGMODE = "NOREG";
    defparam \genblk1.mem1 .RESETMODE = "SYNC";
    defparam \genblk1.mem1 .ASYNC_RESET_RELEASE = "SYNC";
    defparam \genblk1.mem1 .CSDECODE_W = "0b000";
    defparam \genblk1.mem1 .CSDECODE_R = "0b000";
    defparam \genblk1.mem1 .INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem1 .INIT_DATA = "STATIC";
    LUT4 n40157_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6914), .D(n40157), 
         .Z(n40158)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40157_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40152_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6916), .D(n40152), 
         .Z(n40153)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40152_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40147_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6918), .D(n40147), 
         .Z(n40148)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40147_bdd_3_lut_4_lut.init = 16'hf780;
    PDPW16KD \genblk1.mem0  (.DI0(icache_refill_data[0]), .DI1(icache_refill_data[1]), 
            .DI2(icache_refill_data[2]), .DI3(icache_refill_data[3]), .DI4(icache_refill_data[4]), 
            .DI5(icache_refill_data[5]), .DI6(icache_refill_data[6]), .DI7(icache_refill_data[7]), 
            .DI8(icache_refill_data[8]), .DI9(icache_refill_data[9]), .DI10(icache_refill_data[10]), 
            .DI11(icache_refill_data[11]), .DI12(icache_refill_data[12]), 
            .DI13(icache_refill_data[13]), .DI14(icache_refill_data[14]), 
            .DI15(icache_refill_data[15]), .DI16(icache_refill_data[16]), 
            .DI17(icache_refill_data[17]), .DI18(icache_refill_data[18]), 
            .DI19(icache_refill_data[19]), .DI20(icache_refill_data[20]), 
            .DI21(icache_refill_data[21]), .DI22(icache_refill_data[22]), 
            .DI23(icache_refill_data[23]), .DI24(icache_refill_data[24]), 
            .DI25(icache_refill_data[25]), .DI26(icache_refill_data[26]), 
            .DI27(icache_refill_data[27]), .DI28(icache_refill_data[28]), 
            .DI29(icache_refill_data[29]), .DI30(icache_refill_data[30]), 
            .DI31(icache_refill_data[31]), .DI32(GND_net), .DI33(GND_net), 
            .DI34(GND_net), .DI35(GND_net), .ADW0(\dmem_write_address[0] ), 
            .ADW1(\dmem_write_address[1] ), .ADW2(\icache_refill_address[4] ), 
            .ADW3(\icache_refill_address[5] ), .ADW4(\icache_refill_address[6] ), 
            .ADW5(\icache_refill_address[7] ), .ADW6(\icache_refill_address[8] ), 
            .ADW7(\icache_refill_address[9] ), .ADW8(\icache_refill_address[10] ), 
            .BE0(VCC_net), .BE1(VCC_net), .BE2(VCC_net), .BE3(VCC_net), 
            .CEW(REF_CLK_c_enable_44), .CLKW(REF_CLK_c), .CSW0(GND_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(GND_net), .ADR5(n6837[0]), 
            .ADR6(n6837[1]), .ADR7(n6837[2]), .ADR8(n6837[3]), .ADR9(n6837[4]), 
            .ADR10(n6837[5]), .ADR11(n6837[6]), .ADR12(n6837[7]), .ADR13(n6837[8]), 
            .CER(VCC_net), .OCER(VCC_net), .CLKR(REF_CLK_c), .CSR0(GND_net), 
            .CSR1(GND_net), .CSR2(GND_net), .RST(GND_net), .DO0(n7052), 
            .DO1(n7053), .DO2(n7054), .DO3(n7055), .DO4(n7056), .DO5(n7057), 
            .DO6(n7058), .DO7(n7059), .DO8(n7060), .DO9(n7061), .DO10(n7062), 
            .DO11(n7063), .DO12(n7064), .DO13(n7065), .DO18(n7034), 
            .DO19(n7035), .DO20(n7036), .DO21(n7037), .DO22(n7038), 
            .DO23(n7039), .DO24(n7040), .DO25(n7041), .DO26(n7042), 
            .DO27(n7043), .DO28(n7044), .DO29(n7045), .DO30(n7046), 
            .DO31(n7047), .DO32(n7048), .DO33(n7049), .DO34(n7050), 
            .DO35(n7051));
    defparam \genblk1.mem0 .DATA_WIDTH_W = 36;
    defparam \genblk1.mem0 .DATA_WIDTH_R = 36;
    defparam \genblk1.mem0 .GSR = "DISABLED";
    defparam \genblk1.mem0 .REGMODE = "NOREG";
    defparam \genblk1.mem0 .RESETMODE = "SYNC";
    defparam \genblk1.mem0 .ASYNC_RESET_RELEASE = "SYNC";
    defparam \genblk1.mem0 .CSDECODE_W = "0b000";
    defparam \genblk1.mem0 .CSDECODE_R = "0b000";
    defparam \genblk1.mem0 .INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.mem0 .INIT_DATA = "STATIC";
    FD1S3AX \genblk1.mem  (.D(icache_refill_data[31]), .CK(REF_CLK_c), .Q(n6938));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem .GSR = "ENABLED";
    LUT4 n40139_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6920), .D(n40139), 
         .Z(n40140)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40139_bdd_3_lut_4_lut.init = 16'hf780;
    FD1S3AX \genblk1.mem_2929  (.D(icache_refill_data[30]), .CK(REF_CLK_c), 
            .Q(n6936));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2929 .GSR = "ENABLED";
    LUT4 n40134_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6922), .D(n40134), 
         .Z(n40135)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40134_bdd_3_lut_4_lut.init = 16'hf780;
    FD1S3AX \genblk1.mem_2928  (.D(icache_refill_data[29]), .CK(REF_CLK_c), 
            .Q(n6934));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2928 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2927  (.D(icache_refill_data[28]), .CK(REF_CLK_c), 
            .Q(n6932));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2927 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2926  (.D(icache_refill_data[27]), .CK(REF_CLK_c), 
            .Q(n6930));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2926 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2925  (.D(icache_refill_data[26]), .CK(REF_CLK_c), 
            .Q(n6928));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2925 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2924  (.D(icache_refill_data[25]), .CK(REF_CLK_c), 
            .Q(n6926));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2924 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2923  (.D(icache_refill_data[24]), .CK(REF_CLK_c), 
            .Q(n6924));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2923 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2922  (.D(icache_refill_data[23]), .CK(REF_CLK_c), 
            .Q(n6922));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2922 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2921  (.D(icache_refill_data[22]), .CK(REF_CLK_c), 
            .Q(n6920));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2921 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2920  (.D(icache_refill_data[21]), .CK(REF_CLK_c), 
            .Q(n6918));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2920 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2919  (.D(icache_refill_data[20]), .CK(REF_CLK_c), 
            .Q(n6916));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2919 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2918  (.D(icache_refill_data[19]), .CK(REF_CLK_c), 
            .Q(n6914));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2918 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2917  (.D(icache_refill_data[18]), .CK(REF_CLK_c), 
            .Q(n6912));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2917 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2916  (.D(icache_refill_data[17]), .CK(REF_CLK_c), 
            .Q(n6910));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2916 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2915  (.D(icache_refill_data[16]), .CK(REF_CLK_c), 
            .Q(n6908));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2915 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2914  (.D(icache_refill_data[15]), .CK(REF_CLK_c), 
            .Q(n6906));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2914 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2913  (.D(icache_refill_data[14]), .CK(REF_CLK_c), 
            .Q(n6904));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2913 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2912  (.D(icache_refill_data[13]), .CK(REF_CLK_c), 
            .Q(n6902));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2912 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2911  (.D(icache_refill_data[12]), .CK(REF_CLK_c), 
            .Q(n6900));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2911 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2910  (.D(icache_refill_data[11]), .CK(REF_CLK_c), 
            .Q(n6898));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2910 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2909  (.D(icache_refill_data[10]), .CK(REF_CLK_c), 
            .Q(n6896));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2909 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2908  (.D(icache_refill_data[9]), .CK(REF_CLK_c), 
            .Q(n6894));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2908 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2907  (.D(icache_refill_data[8]), .CK(REF_CLK_c), 
            .Q(n6892));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2907 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2906  (.D(icache_refill_data[7]), .CK(REF_CLK_c), 
            .Q(n6890));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2906 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2905  (.D(icache_refill_data[6]), .CK(REF_CLK_c), 
            .Q(n6888));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2905 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2904  (.D(icache_refill_data[5]), .CK(REF_CLK_c), 
            .Q(n6886));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2904 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2903  (.D(icache_refill_data[4]), .CK(REF_CLK_c), 
            .Q(n6884));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2903 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2902  (.D(icache_refill_data[3]), .CK(REF_CLK_c), 
            .Q(n6882));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2902 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2901  (.D(icache_refill_data[2]), .CK(REF_CLK_c), 
            .Q(n6880));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2901 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2900  (.D(icache_refill_data[1]), .CK(REF_CLK_c), 
            .Q(n6878));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2900 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2899  (.D(icache_refill_data[0]), .CK(REF_CLK_c), 
            .Q(n6876));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(291[26:33])
    defparam \genblk1.mem_2899 .GSR = "ENABLED";
    LUT4 n40129_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6924), .D(n40129), 
         .Z(n40130)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40129_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40124_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6926), .D(n40124), 
         .Z(n40125)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40124_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40119_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6928), .D(n40119), 
         .Z(n40120)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40119_bdd_3_lut_4_lut.init = 16'hf780;
    FD1S3AX \genblk1.mem_2898  (.D(icache_refill_ready), .CK(REF_CLK_c), 
            .Q(n6873));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2898 .GSR = "ENABLED";
    LUT4 n40114_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6930), .D(n40114), 
         .Z(n40115)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40114_bdd_3_lut_4_lut.init = 16'hf780;
    FD1S3AX \genblk1.mem_2894  (.D(\icache_refill_address[12] ), .CK(REF_CLK_c), 
            .Q(n6870));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_2894 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2892  (.D(\icache_refill_address[11] ), .CK(REF_CLK_c), 
            .Q(n6868));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_2892 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2891  (.D(n6837[8]), .CK(REF_CLK_c), .Q(\genblk1.ra [8]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2891 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2890  (.D(\icache_refill_address[10] ), .CK(REF_CLK_c), 
            .Q(n6866));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_2890 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2889  (.D(n6837[7]), .CK(REF_CLK_c), .Q(\genblk1.ra [7]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2889 .GSR = "ENABLED";
    LUT4 n40109_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6932), .D(n40109), 
         .Z(n40110)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40109_bdd_3_lut_4_lut.init = 16'hf780;
    FD1S3AX \genblk1.mem_2888  (.D(\icache_refill_address[9] ), .CK(REF_CLK_c), 
            .Q(n6864));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_2888 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2887  (.D(n6837[6]), .CK(REF_CLK_c), .Q(\genblk1.ra [6]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2887 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2886  (.D(\icache_refill_address[8] ), .CK(REF_CLK_c), 
            .Q(n6862));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_2886 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2885  (.D(n6837[5]), .CK(REF_CLK_c), .Q(\genblk1.ra [5]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2885 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2884  (.D(\icache_refill_address[7] ), .CK(REF_CLK_c), 
            .Q(n6860));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_2884 .GSR = "ENABLED";
    LUT4 n40104_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6934), .D(n40104), 
         .Z(n40105)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40104_bdd_3_lut_4_lut.init = 16'hf780;
    FD1S3AX \genblk1.mem_2883  (.D(n6837[4]), .CK(REF_CLK_c), .Q(\genblk1.ra [4]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2883 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2882  (.D(\icache_refill_address[6] ), .CK(REF_CLK_c), 
            .Q(n6858));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_2882 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2881  (.D(n6837[3]), .CK(REF_CLK_c), .Q(\genblk1.ra [3]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2881 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2880  (.D(\icache_refill_address[5] ), .CK(REF_CLK_c), 
            .Q(n6856));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_2880 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2879  (.D(n6837[2]), .CK(REF_CLK_c), .Q(\genblk1.ra [2]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2879 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2878  (.D(\icache_refill_address[4] ), .CK(REF_CLK_c), 
            .Q(n6854));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_2878 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2877  (.D(n6837[1]), .CK(REF_CLK_c), .Q(\genblk1.ra [1]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2877 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2876  (.D(\dmem_write_address[1] ), .CK(REF_CLK_c), 
            .Q(n6852));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_2876 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2875  (.D(n6837[0]), .CK(REF_CLK_c), .Q(\genblk1.ra [0]));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.mem_2875 .GSR = "ENABLED";
    FD1S3AX \genblk1.mem_2874  (.D(\dmem_write_address[0] ), .CK(REF_CLK_c), 
            .Q(n6850));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam \genblk1.mem_2874 .GSR = "ENABLED";
    LUT4 n40096_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6936), .D(n40096), 
         .Z(n40097)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40096_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40091_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6938), .D(n40091), 
         .Z(n40092)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40091_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40269_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6876), .D(n40269), 
         .Z(n40270)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40269_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40070_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6898), .D(n40070), 
         .Z(n40071)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40070_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 i31976_2_lut_3_lut (.A(n6873), .B(n6872), .C(\genblk1.ra[10] ), 
         .Z(n37144)) /* synthesis lut_function=(!(A (B+(C))+!A (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam i31976_2_lut_3_lut.init = 16'h0707;
    LUT4 n40075_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6900), .D(n40075), 
         .Z(n40076)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40075_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40279_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6904), .D(n40279), 
         .Z(n40280)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40279_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_2872_i1_3_lut (.A(\pc_a[2] ), .B(\genblk1.ra [0]), .C(n45183), 
         .Z(n6837[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_2872_i1_3_lut.init = 16'hcaca;
    LUT4 mux_2872_i2_3_lut (.A(\pc_a[3] ), .B(\genblk1.ra [1]), .C(n45183), 
         .Z(n6837[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_2872_i2_3_lut.init = 16'hcaca;
    CCU2C equal_2894_9 (.A0(\genblk1.ra [7]), .B0(n6864), .C0(\genblk1.ra [6]), 
          .D0(n6862), .A1(\genblk1.ra [5]), .B1(n6860), .C1(\genblk1.ra [4]), 
          .D1(n6858), .CIN(n27352), .COUT(n27353));
    defparam equal_2894_9.INIT0 = 16'h9009;
    defparam equal_2894_9.INIT1 = 16'h9009;
    defparam equal_2894_9.INJECT1_0 = "YES";
    defparam equal_2894_9.INJECT1_1 = "YES";
    LUT4 mux_2872_i3_3_lut (.A(\pc_a[4] ), .B(\genblk1.ra [2]), .C(n45183), 
         .Z(n6837[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_2872_i3_3_lut.init = 16'hcaca;
    LUT4 mux_2872_i4_3_lut (.A(\pc_a[5] ), .B(\genblk1.ra [3]), .C(n45183), 
         .Z(n6837[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_2872_i4_3_lut.init = 16'hcaca;
    LUT4 mux_2872_i5_3_lut (.A(\pc_a[6] ), .B(\genblk1.ra [4]), .C(n45183), 
         .Z(n6837[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_2872_i5_3_lut.init = 16'hcaca;
    LUT4 mux_2872_i6_3_lut (.A(\pc_a[7] ), .B(\genblk1.ra [5]), .C(n45183), 
         .Z(n6837[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_2872_i6_3_lut.init = 16'hcaca;
    LUT4 mux_2872_i7_3_lut (.A(\pc_a[8] ), .B(\genblk1.ra [6]), .C(n45183), 
         .Z(n6837[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_2872_i7_3_lut.init = 16'hcaca;
    LUT4 mux_2872_i8_3_lut (.A(\pc_a[9] ), .B(\genblk1.ra [7]), .C(n45183), 
         .Z(n6837[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_2872_i8_3_lut.init = 16'hcaca;
    LUT4 mux_2872_i9_3_lut (.A(\pc_a[10] ), .B(\genblk1.ra [8]), .C(n45183), 
         .Z(n6837[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam mux_2872_i9_3_lut.init = 16'hcaca;
    FD1P3AX \genblk1.ra_rep_8__0_i0  (.D(\pc_a[11] ), .SP(REF_CLK_c_enable_1178), 
            .CK(REF_CLK_c), .Q(\genblk1.ra[9] ));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.ra_rep_8__0_i0 .GSR = "ENABLED";
    CCU2C equal_2894_0 (.A0(\genblk1.ra[10] ), .B0(n6870), .C0(GND_net), 
          .D0(VCC_net), .A1(\genblk1.ra[9] ), .B1(n6868), .C1(\genblk1.ra [8]), 
          .D1(n6866), .COUT(n27352));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam equal_2894_0.INIT0 = 16'h0009;
    defparam equal_2894_0.INIT1 = 16'h9009;
    defparam equal_2894_0.INJECT1_0 = "NO";
    defparam equal_2894_0.INJECT1_1 = "YES";
    CCU2C equal_2894_11 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n27354), 
          .S0(n6872));
    defparam equal_2894_11.INIT0 = 16'h0000;
    defparam equal_2894_11.INIT1 = 16'h0000;
    defparam equal_2894_11.INJECT1_0 = "NO";
    defparam equal_2894_11.INJECT1_1 = "NO";
    CCU2C equal_2894_11_22475 (.A0(\genblk1.ra [3]), .B0(n6856), .C0(\genblk1.ra [2]), 
          .D0(n6854), .A1(\genblk1.ra [1]), .B1(n6852), .C1(\genblk1.ra [0]), 
          .D1(n6850), .CIN(n27353), .COUT(n27354));
    defparam equal_2894_11_22475.INIT0 = 16'h9009;
    defparam equal_2894_11_22475.INIT1 = 16'h9009;
    defparam equal_2894_11_22475.INJECT1_0 = "YES";
    defparam equal_2894_11_22475.INJECT1_1 = "YES";
    FD1P3AX \genblk1.ra_i10  (.D(\pc_a[12] ), .SP(REF_CLK_c_enable_1425), 
            .CK(REF_CLK_c), .Q(\genblk1.ra[10] ));   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam \genblk1.ra_i10 .GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut (.A(icache_refill_ready), .B(\icache_refill_address[11] ), 
         .C(\icache_refill_address[12] ), .Z(REF_CLK_c_enable_43)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_360 (.A(icache_refill_ready), .B(\icache_refill_address[11] ), 
         .C(\icache_refill_address[12] ), .Z(REF_CLK_c_enable_44)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam i1_2_lut_3_lut_adj_360.init = 16'h0202;
    LUT4 i1_2_lut_3_lut_adj_361 (.A(icache_refill_ready), .B(\icache_refill_address[11] ), 
         .C(\icache_refill_address[12] ), .Z(REF_CLK_c_enable_36)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam i1_2_lut_3_lut_adj_361.init = 16'h0808;
    LUT4 i1_2_lut_3_lut_adj_362 (.A(icache_refill_ready), .B(\icache_refill_address[11] ), 
         .C(\icache_refill_address[12] ), .Z(REF_CLK_c_enable_42)) /* synthesis lut_function=(A (B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(299[4:22])
    defparam i1_2_lut_3_lut_adj_362.init = 16'h8080;
    LUT4 n40236_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6902), .D(n40236), 
         .Z(n40237)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40236_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40230_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6878), .D(n40230), 
         .Z(n40231)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40230_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40225_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6880), .D(n40225), 
         .Z(n40226)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40225_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40220_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6882), .D(n40220), 
         .Z(n40221)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40220_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40212_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6884), .D(n40212), 
         .Z(n40213)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40212_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40207_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6886), .D(n40207), 
         .Z(n40208)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40207_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40202_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6888), .D(n40202), 
         .Z(n40203)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40202_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40197_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6890), .D(n40197), 
         .Z(n40198)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40197_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40192_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6892), .D(n40192), 
         .Z(n40193)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40192_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40187_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6894), .D(n40187), 
         .Z(n40188)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40187_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40182_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6896), .D(n40182), 
         .Z(n40183)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40182_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40177_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6906), .D(n40177), 
         .Z(n40178)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40177_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40172_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6908), .D(n40172), 
         .Z(n40173)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40172_bdd_3_lut_4_lut.init = 16'hf780;
    LUT4 n40167_bdd_3_lut_4_lut (.A(n6873), .B(n6872), .C(n6910), .D(n40167), 
         .Z(n40168)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_ram.v(302[14] 304[26])
    defparam n40167_bdd_3_lut_4_lut.init = 16'hf780;
    
endmodule
//
// Verilog Description of module \lm32_debug(watchpoints=32'b0) 
//

module \lm32_debug(watchpoints=32'b0)  (dc_re, REF_CLK_c, REF_CLK_c_enable_388, 
            REF_CLK_c_enable_1606, n36336) /* synthesis syn_module_defined=1 */ ;
    output dc_re;
    input REF_CLK_c;
    input REF_CLK_c_enable_388;
    input REF_CLK_c_enable_1606;
    input n36336;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    
    FD1P3DX dc_re_10 (.D(n36336), .SP(REF_CLK_c_enable_388), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(dc_re)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=1216, LSE_RLINE=1249 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_debug.v(296[5] 299[8])
    defparam dc_re_10.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module lm32_decoder
//

module lm32_decoder (n45106, n41365, n41362, n11807, n41244, n41247, 
            n6028, n41295, n45075, VCC_net, n6777, n11834, n41228, 
            n20863, n41198, n30058, n41381, \bypass_data_0[0] , \d_result_0[0] , 
            \bypass_data_0[1] , \d_result_0[1] , n41363, n31717, bret_d, 
            n6779, \genblk1.wait_one_tick_done , n6780, n6770, n6781, 
            n6775, n6776, n10475, n41382, n6778, eret_d, n41364, 
            n41285, load_d, n32910, n32356, n10, store_d, n41361, 
            break_d, n41367, valid_d, n10_adj_145, n30070, n41196, 
            n30888, n41291, n41373, n41208, n31207, \instruction_d[13] , 
            n31218, \instruction_d[12] , n31219, n31542, branch_d, 
            write_enable_d, n41227, n41229, n41281, \instruction_d[11] , 
            n31221, n41377, n31216, n41376, n31212, n41375, n31220, 
            n31213, n41368, n31217, n41374, n31214, n41371, n31211, 
            n41372, n31209, n41348, n31206, n41370, n31210, n41369, 
            n31215, \instruction_d[14] , n31208, branch_predict_taken_d, 
            n41179, n30820, n41175, adder_op_d_N_1366, n6026, n41187, 
            valid_f, n41203, n31132, n45181, valid_f_N_1250, bypass_data_1, 
            n31309, n31310, n31323, n31298, n31300, n31322, n31302, 
            n31316, n31304, \extended_immediate[31] , n31320, n31317, 
            n41452, n31306, n31295, n31311, n31313, n31315, n31319, 
            n31321, n31296, n31314, n31318, n31308, n31294, n31325, 
            n31312, n31324, n31297, n31299, n31301, n31303, n31305, 
            n31307, x_bypass_enable_d, x_result_sel_csr_d, n41296, n41248, 
            n41441, n41319, n45105, n41241, n30216, n31519, m_bypass_enable_d, 
            n41408, n6760, n2, n19987, n31549, n6761, n2_adj_146, 
            n6762, n2_adj_147, n6763, n2_adj_148, m_result_sel_compare_d, 
            n41451, n6768, n6764, n10589, n45183, n40093, n40094, 
            n6766, n10585, n6769, n10591, n41419, n10485, x_bypass_enable_x, 
            n32006, m_bypass_enable_m, n31984, n10593, n6767, n10587, 
            n41312, n41437, n41184, n37939, n41366, n41201, \d_result_sel_1_d[1] , 
            n6771, n10595, n37933, n41205, n37934, n37936, n6765, 
            n10452, n37937, n37938, n37935, n31494) /* synthesis syn_module_defined=1 */ ;
    input n45106;
    input n41365;
    input n41362;
    output n11807;
    output n41244;
    input n41247;
    input n6028;
    input n41295;
    output n45075;
    input VCC_net;
    input n6777;
    output n11834;
    input n41228;
    output n20863;
    output n41198;
    output n30058;
    input n41381;
    input \bypass_data_0[0] ;
    output \d_result_0[0] ;
    input \bypass_data_0[1] ;
    output \d_result_0[1] ;
    input n41363;
    input n31717;
    output bret_d;
    input n6779;
    input \genblk1.wait_one_tick_done ;
    input n6780;
    input n6770;
    input n6781;
    input n6775;
    input n6776;
    output n10475;
    input n41382;
    input n6778;
    output eret_d;
    output n41364;
    input n41285;
    output load_d;
    output n32910;
    output n32356;
    input n10;
    output store_d;
    input n41361;
    output break_d;
    input n41367;
    input valid_d;
    output n10_adj_145;
    input n30070;
    output n41196;
    input n30888;
    output n41291;
    input n41373;
    input n41208;
    output n31207;
    input \instruction_d[13] ;
    output n31218;
    input \instruction_d[12] ;
    output n31219;
    input n31542;
    output branch_d;
    output write_enable_d;
    input n41227;
    input n41229;
    input n41281;
    input \instruction_d[11] ;
    output n31221;
    input n41377;
    output n31216;
    input n41376;
    output n31212;
    input n41375;
    output n31220;
    output n31213;
    input n41368;
    output n31217;
    input n41374;
    output n31214;
    input n41371;
    output n31211;
    input n41372;
    output n31209;
    input n41348;
    output n31206;
    input n41370;
    output n31210;
    input n41369;
    output n31215;
    input \instruction_d[14] ;
    output n31208;
    output branch_predict_taken_d;
    output n41179;
    input n30820;
    output n41175;
    output adder_op_d_N_1366;
    output n6026;
    output n41187;
    input valid_f;
    input n41203;
    output n31132;
    input n45181;
    output valid_f_N_1250;
    input [31:0]bypass_data_1;
    output n31309;
    output n31310;
    output n31323;
    output n31298;
    output n31300;
    output n31322;
    output n31302;
    output n31316;
    output n31304;
    output \extended_immediate[31] ;
    output n31320;
    output n31317;
    input n41452;
    output n31306;
    output n31295;
    output n31311;
    output n31313;
    output n31315;
    output n31319;
    output n31321;
    output n31296;
    output n31314;
    output n31318;
    output n31308;
    output n31294;
    output n31325;
    output n31312;
    output n31324;
    output n31297;
    output n31299;
    output n31301;
    output n31303;
    output n31305;
    output n31307;
    output x_bypass_enable_d;
    output x_result_sel_csr_d;
    input n41296;
    input n41248;
    output n41441;
    output n41319;
    input n45105;
    input n41241;
    input n30216;
    input n31519;
    output m_bypass_enable_d;
    output n41408;
    input n6760;
    output n2;
    input n19987;
    output n31549;
    input n6761;
    output n2_adj_146;
    input n6762;
    output n2_adj_147;
    input n6763;
    output n2_adj_148;
    output m_result_sel_compare_d;
    output n41451;
    input n6768;
    input n6764;
    output n10589;
    input n45183;
    input n40093;
    output n40094;
    input n6766;
    output n10585;
    input n6769;
    output n10591;
    output n41419;
    output n10485;
    input x_bypass_enable_x;
    output n32006;
    input m_bypass_enable_m;
    output n31984;
    output n10593;
    input n6767;
    output n10587;
    output n41312;
    input n41437;
    output n41184;
    output n37939;
    input n41366;
    output n41201;
    output \d_result_sel_1_d[1] ;
    input n6771;
    output n10595;
    output n37933;
    output n41205;
    output n37934;
    output n37936;
    input n6765;
    output n10452;
    output n37937;
    output n37938;
    output n37935;
    output n31494;
    
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    
    wire n41438, n31427, n34908, n34760, n41462, n27797, n41287, 
        n41214, n11849, n32522, n32516, n32512, n35068, n30184, 
        n30904, n10479, n41294, n35012, n35086, n41286, n41188, 
        n41192, n41204, n11815, n35016, n41280, n45069, n10487, 
        n41440, n34474, n29801, n45070, n10473, n41206, n31505, 
        n42801, n41213, n34912, n30136, n34766, n31675, n19888, 
        n41439, n33940, n34578, n34570, n31829;
    
    LUT4 i1_3_lut_4_lut (.A(n45106), .B(n41438), .C(n41365), .D(n41362), 
         .Z(n11807)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_3_lut_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n41244), .B(n41247), .C(n6028), .D(n31427), 
         .Z(n34908)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(376[20:65])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0e00;
    LUT4 i1_2_lut_4_lut_4_lut (.A(n41244), .B(n41247), .C(n41295), .D(n45075), 
         .Z(n34760)) /* synthesis lut_function=(!(A+(B ((D)+!C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(376[20:65])
    defparam i1_2_lut_4_lut_4_lut.init = 16'h1151;
    PFUMX i34361 (.BLUT(n41462), .ALUT(VCC_net), .C0(n6777), .Z(n27797));
    LUT4 i15577_2_lut_3_lut_4_lut (.A(n41287), .B(n11834), .C(n11807), 
         .D(n41228), .Z(n20863)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(348[20:68])
    defparam i15577_2_lut_3_lut_4_lut.init = 16'heee0;
    LUT4 i33097_3_lut_rep_793_4_lut (.A(n31427), .B(n41214), .C(n11849), 
         .D(n27797), .Z(n41198)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i33097_3_lut_rep_793_4_lut.init = 16'h0800;
    LUT4 i14575_2_lut_4_lut (.A(n41295), .B(n30058), .C(n41381), .D(\bypass_data_0[0] ), 
         .Z(\d_result_0[0] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(D))) */ ;
    defparam i14575_2_lut_4_lut.init = 16'h7f00;
    LUT4 i15000_2_lut_4_lut (.A(n41295), .B(n30058), .C(n41381), .D(\bypass_data_0[1] ), 
         .Z(\d_result_0[1] )) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(D))) */ ;
    defparam i15000_2_lut_4_lut.init = 16'h7f00;
    LUT4 i33163_4_lut (.A(n41363), .B(n41365), .C(n31717), .D(n32522), 
         .Z(bret_d)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(346[20:67])
    defparam i33163_4_lut.init = 16'h0010;
    LUT4 i1_4_lut (.A(n6779), .B(\genblk1.wait_one_tick_done ), .C(n6780), 
         .D(n32516), .Z(n32522)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_4_lut.init = 16'hff7f;
    LUT4 i1_2_lut (.A(n6770), .B(n6781), .Z(n32516)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut.init = 16'hdddd;
    LUT4 i5134_2_lut (.A(n6775), .B(n6776), .Z(n10475)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(359[20:68])
    defparam i5134_2_lut.init = 16'heeee;
    LUT4 i33166_4_lut (.A(n41382), .B(n32512), .C(n6770), .D(n6778), 
         .Z(eret_d)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(346[20:67])
    defparam i33166_4_lut.init = 16'h1113;
    LUT4 i1_3_lut (.A(n41363), .B(n31717), .C(n41364), .Z(n32512)) /* synthesis lut_function=(A+((C)+!B)) */ ;
    defparam i1_3_lut.init = 16'hfbfb;
    LUT4 i33183_4_lut (.A(n35068), .B(n30184), .C(n30904), .D(n41285), 
         .Z(load_d)) /* synthesis lut_function=(!(A (B (C))+!A (B (C (D))))) */ ;
    defparam i33183_4_lut.init = 16'h3f7f;
    LUT4 i1_4_lut_adj_279 (.A(n41382), .B(n41363), .C(n32910), .D(n32356), 
         .Z(n30904)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;
    defparam i1_4_lut_adj_279.init = 16'hffec;
    LUT4 i5137_2_lut (.A(n6779), .B(n6780), .Z(n10479)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(367[20:68])
    defparam i5137_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_280 (.A(n6778), .B(n6780), .Z(n32910)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(367[20:68])
    defparam i1_2_lut_adj_280.init = 16'heeee;
    LUT4 i33178_3_lut_4_lut (.A(n41294), .B(n41285), .C(n10), .D(n35012), 
         .Z(store_d)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B (C (D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(349[20:68])
    defparam i33178_3_lut_4_lut.init = 16'h01ff;
    LUT4 i33095_3_lut_4_lut (.A(n41294), .B(n41285), .C(n35086), .D(n41361), 
         .Z(break_d)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(349[20:68])
    defparam i33095_3_lut_4_lut.init = 16'h0001;
    LUT4 i3_2_lut_3_lut_4_lut (.A(n41367), .B(n41286), .C(valid_d), .D(n41287), 
         .Z(n10_adj_145)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(353[20:69])
    defparam i3_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_791_3_lut_4_lut (.A(n41367), .B(n41286), .C(n30070), 
         .D(n41287), .Z(n41196)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(353[20:69])
    defparam i1_2_lut_rep_791_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_3_lut_4_lut_adj_281 (.A(n41367), .B(n41286), .C(n30888), .D(n10), 
         .Z(n30184)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(353[20:69])
    defparam i1_3_lut_4_lut_adj_281.init = 16'hff0e;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n41291), .B(n41373), .C(n41208), .D(n41188), 
         .Z(n31207)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'h0444;
    LUT4 i1_3_lut_4_lut_4_lut_adj_282 (.A(n41291), .B(\instruction_d[13] ), 
         .C(n41208), .D(n41188), .Z(n31218)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_282.init = 16'h0444;
    LUT4 i1_3_lut_4_lut_4_lut_adj_283 (.A(n41291), .B(\instruction_d[12] ), 
         .C(n41208), .D(n41188), .Z(n31219)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_283.init = 16'h0444;
    LUT4 i33174_4_lut (.A(n41192), .B(n41204), .C(n41287), .D(n31542), 
         .Z(branch_d)) /* synthesis lut_function=(!(A (B+!((D)+!C)))) */ ;
    defparam i33174_4_lut.init = 16'h7757;
    LUT4 i1_4_lut_adj_284 (.A(n41192), .B(store_d), .C(n11815), .D(n35016), 
         .Z(write_enable_d)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_4_lut_adj_284.init = 16'h2000;
    LUT4 i1_4_lut_adj_285 (.A(n35068), .B(n41227), .C(n41229), .D(n41281), 
         .Z(n35012)) /* synthesis lut_function=(A (B+(D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_285.init = 16'hfac8;
    LUT4 i1_3_lut_4_lut_4_lut_adj_286 (.A(n41291), .B(\instruction_d[11] ), 
         .C(n41208), .D(n41188), .Z(n31221)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_286.init = 16'h0444;
    LUT4 i1_3_lut_4_lut_4_lut_adj_287 (.A(n41291), .B(n41377), .C(n41208), 
         .D(n41188), .Z(n31216)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_287.init = 16'h0444;
    LUT4 i1_3_lut_4_lut_4_lut_adj_288 (.A(n41291), .B(n41376), .C(n41208), 
         .D(n41188), .Z(n31212)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_288.init = 16'h0444;
    LUT4 i1_3_lut_4_lut_4_lut_adj_289 (.A(n41291), .B(n41375), .C(n41208), 
         .D(n41188), .Z(n31220)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_289.init = 16'h0444;
    LUT4 i1_3_lut_4_lut_4_lut_adj_290 (.A(n41291), .B(n41361), .C(n41208), 
         .D(n41188), .Z(n31213)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_290.init = 16'h0444;
    LUT4 i1_3_lut_4_lut_4_lut_adj_291 (.A(n41291), .B(n41368), .C(n41208), 
         .D(n41188), .Z(n31217)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_291.init = 16'h0444;
    LUT4 i1_3_lut_4_lut_4_lut_adj_292 (.A(n41291), .B(n41374), .C(n41208), 
         .D(n41188), .Z(n31214)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_292.init = 16'h0444;
    LUT4 i1_3_lut_4_lut_4_lut_adj_293 (.A(n41291), .B(n41371), .C(n41208), 
         .D(n41188), .Z(n31211)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_293.init = 16'h0444;
    LUT4 i1_3_lut_4_lut_4_lut_adj_294 (.A(n41291), .B(n41372), .C(n41208), 
         .D(n41188), .Z(n31209)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_294.init = 16'h0444;
    LUT4 i1_3_lut_4_lut_4_lut_adj_295 (.A(n41291), .B(n41348), .C(n41208), 
         .D(n41188), .Z(n31206)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_295.init = 16'h0444;
    LUT4 i1_3_lut_4_lut_4_lut_adj_296 (.A(n41291), .B(n41370), .C(n41208), 
         .D(n41188), .Z(n31210)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_296.init = 16'h0444;
    LUT4 i1_3_lut_4_lut_4_lut_adj_297 (.A(n41291), .B(n41369), .C(n41208), 
         .D(n41188), .Z(n31215)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_297.init = 16'h0444;
    LUT4 i1_3_lut_4_lut_4_lut_adj_298 (.A(n41291), .B(\instruction_d[14] ), 
         .C(n41208), .D(n41188), .Z(n31208)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_298.init = 16'h0444;
    LUT4 i1_4_lut_adj_299 (.A(n41281), .B(n41280), .C(n45069), .D(n41348), 
         .Z(branch_predict_taken_d)) /* synthesis lut_function=(!(A (B)+!A (B (C+!(D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(414[8:26])
    defparam i1_4_lut_adj_299.init = 16'h3733;
    LUT4 i5145_2_lut (.A(n6776), .B(n6777), .Z(n10487)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(346[20:67])
    defparam i5145_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_rep_875_4_lut (.A(n10475), .B(n41382), .C(n6777), .D(n31542), 
         .Z(n41280)) /* synthesis lut_function=(A (B+!(D))+!A (B (C+!(D))+!B !(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(346[20:67])
    defparam i1_2_lut_rep_875_4_lut.init = 16'hc8ff;
    LUT4 i1_2_lut_rep_882_4_lut (.A(n41440), .B(\genblk1.wait_one_tick_done ), 
         .C(n6780), .D(n41365), .Z(n41287)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i1_2_lut_rep_882_4_lut.init = 16'hffbf;
    LUT4 i15456_2_lut_rep_774_3_lut_4_lut (.A(n41281), .B(n45069), .C(n41208), 
         .D(n34474), .Z(n41179)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B (C)))) */ ;
    defparam i15456_2_lut_rep_774_3_lut_4_lut.init = 16'h0fef;
    LUT4 instruction_30__I_0_171_i7_2_lut_3_lut_4_lut_4_lut_rep_1055 (.A(\genblk1.wait_one_tick_done ), 
         .B(n6778), .C(n6781), .D(n6779), .Z(n45075)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam instruction_30__I_0_171_i7_2_lut_3_lut_4_lut_4_lut_rep_1055.init = 16'hfff7;
    LUT4 i1_3_lut_rep_770_4_lut (.A(n41280), .B(n41192), .C(n30820), .D(n29801), 
         .Z(n41175)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_3_lut_rep_770_4_lut.init = 16'hff7f;
    LUT4 i38_1_lut_3_lut_4_lut (.A(n41280), .B(n41192), .C(n30820), .D(n29801), 
         .Z(adder_op_d_N_1366)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i38_1_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_783_3_lut_4_lut (.A(n45070), .B(n41229), .C(n34474), 
         .D(n41281), .Z(n41188)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C+!(D))) */ ;
    defparam i1_2_lut_rep_783_3_lut_4_lut.init = 16'hf0f7;
    LUT4 i2_4_lut (.A(n30058), .B(n41382), .C(n6778), .D(n10473), .Z(n6026)) /* synthesis lut_function=(!((B (C+(D)))+!A)) */ ;
    defparam i2_4_lut.init = 16'h222a;
    LUT4 i5132_2_lut (.A(n6776), .B(n6777), .Z(n10473)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5132_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_rep_782 (.A(branch_predict_taken_d), .B(valid_d), .Z(n41187)) /* synthesis lut_function=(A (B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(414[8:26])
    defparam i1_2_lut_rep_782.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_300 (.A(branch_predict_taken_d), .B(valid_d), 
         .C(valid_f), .D(n41203), .Z(n31132)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(414[8:26])
    defparam i1_3_lut_4_lut_adj_300.init = 16'h0070;
    LUT4 i1_3_lut_4_lut_adj_301 (.A(branch_predict_taken_d), .B(valid_d), 
         .C(n41203), .D(n45181), .Z(valid_f_N_1250)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/spi/rtl/verilog/wb_spi.v(414[8:26])
    defparam i1_3_lut_4_lut_adj_301.init = 16'hfff8;
    LUT4 i1_2_lut_3_lut_4_lut_adj_302 (.A(n34474), .B(n41192), .C(bypass_data_1[0]), 
         .D(n41208), .Z(n31309)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_302.init = 16'hb000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_303 (.A(n34474), .B(n41192), .C(bypass_data_1[2]), 
         .D(n41208), .Z(n31310)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_303.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_304 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[14]), 
         .Z(n31323)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_304.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_305 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[13]), 
         .Z(n31298)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_305.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_306 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[12]), 
         .Z(n31300)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_306.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_307 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[11]), 
         .Z(n31322)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_307.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_308 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[10]), 
         .Z(n31302)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_308.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_309 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[9]), 
         .Z(n31316)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_309.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_310 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[8]), 
         .Z(n31304)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_310.init = 16'hb000;
    LUT4 sign_extend_immediate_I_0_2_lut_4_lut (.A(n41206), .B(n27797), 
         .C(n11849), .D(n41348), .Z(\extended_immediate[31] )) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(586[32:100])
    defparam sign_extend_immediate_I_0_2_lut_4_lut.init = 16'h0800;
    LUT4 i1_3_lut_4_lut_adj_311 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[24]), 
         .Z(n31320)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_311.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_312 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[23]), 
         .Z(n31317)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_312.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_313 (.A(n41365), .B(n41452), .C(n41295), .D(n31505), 
         .Z(n11849)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_313.init = 16'h0080;
    LUT4 i1_3_lut_4_lut_adj_314 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[22]), 
         .Z(n31306)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_314.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_315 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[21]), 
         .Z(n31295)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_315.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_316 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[20]), 
         .Z(n31311)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_316.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_317 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[19]), 
         .Z(n31313)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_317.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_318 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[18]), 
         .Z(n31315)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_318.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_319 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[17]), 
         .Z(n31319)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_319.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_320 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[16]), 
         .Z(n31321)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_320.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_321 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[15]), 
         .Z(n31296)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_321.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_322 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[7]), 
         .Z(n31314)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_322.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_323 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[6]), 
         .Z(n31318)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_323.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_324 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[5]), 
         .Z(n31308)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_324.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_325 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[4]), 
         .Z(n31294)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_325.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_326 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[3]), 
         .Z(n31325)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_326.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_327 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[1]), 
         .Z(n31312)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_327.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_328 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[31]), 
         .Z(n31324)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_328.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_329 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[30]), 
         .Z(n31297)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_329.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_330 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[29]), 
         .Z(n31299)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_330.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_331 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[28]), 
         .Z(n31301)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_331.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_332 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[27]), 
         .Z(n31303)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_332.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_333 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[26]), 
         .Z(n31305)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_333.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_334 (.A(n34474), .B(n41192), .C(n41208), .D(bypass_data_1[25]), 
         .Z(n31307)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_334.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_335 (.A(n41294), .B(n41367), .C(n10475), .D(n41382), 
         .Z(n31505)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(356[20:66])
    defparam i1_3_lut_4_lut_adj_335.init = 16'he000;
    LUT4 i1_2_lut_rep_801_3_lut_4_lut (.A(n41294), .B(n41367), .C(n31427), 
         .D(n41247), .Z(n41206)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(356[20:66])
    defparam i1_2_lut_rep_801_3_lut_4_lut.init = 16'hf0e0;
    LUT4 n6775_bdd_4_lut_35551 (.A(n6775), .B(n6777), .C(n6776), .D(n6781), 
         .Z(n42801)) /* synthesis lut_function=(A (D)+!A (B+((D)+!C))) */ ;
    defparam n6775_bdd_4_lut_35551.init = 16'hff45;
    LUT4 i1_3_lut_rep_808_4_lut (.A(n41294), .B(n41367), .C(n41295), .D(n45075), 
         .Z(n41213)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(356[20:66])
    defparam i1_3_lut_rep_808_4_lut.init = 16'h0010;
    LUT4 i1_4_lut_adj_336 (.A(n34912), .B(n20863), .C(n30136), .D(n34766), 
         .Z(x_bypass_enable_d)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_4_lut_adj_336.init = 16'hff7f;
    LUT4 i1_4_lut_adj_337 (.A(n31427), .B(x_result_sel_csr_d), .C(n31675), 
         .D(n34760), .Z(n34766)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i1_4_lut_adj_337.init = 16'hffdf;
    LUT4 i1_2_lut_adj_338 (.A(n27797), .B(n19888), .Z(n34912)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_338.init = 16'h8888;
    LUT4 i1_4_lut_adj_339 (.A(n41296), .B(n41204), .C(n41439), .D(n41440), 
         .Z(n30136)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(348[20:68])
    defparam i1_4_lut_adj_339.init = 16'hfffe;
    LUT4 i14624_4_lut (.A(n35086), .B(n30888), .C(n41229), .D(n41287), 
         .Z(n19888)) /* synthesis lut_function=(A ((D)+!B)+!A (B (C (D))+!B (C))) */ ;
    defparam i14624_4_lut.init = 16'hfa32;
    LUT4 i2_rep_113_4_lut (.A(n41248), .B(n41441), .C(n33940), .D(n45075), 
         .Z(n31427)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_rep_113_4_lut.init = 16'hfeee;
    LUT4 instruction_30__I_0_183_i9_2_lut_rep_809_3_lut_4_lut (.A(n41319), 
         .B(n41382), .C(n41367), .D(n41294), .Z(n41214)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(374[20:65])
    defparam instruction_30__I_0_183_i9_2_lut_rep_809_3_lut_4_lut.init = 16'hfff8;
    LUT4 n947_bdd_2_lut_35290_rep_1050 (.A(n42801), .B(n45105), .Z(n45070)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam n947_bdd_2_lut_35290_rep_1050.init = 16'hbbbb;
    LUT4 i1_4_lut_adj_340 (.A(n31675), .B(n41241), .C(n11849), .D(n30216), 
         .Z(n29801)) /* synthesis lut_function=((B (C+(D))+!B (C))+!A) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(402[14:76])
    defparam i1_4_lut_adj_340.init = 16'hfdf5;
    LUT4 i1_4_lut_adj_341 (.A(n34578), .B(n29801), .C(n31519), .D(n20863), 
         .Z(m_bypass_enable_d)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(402[14:76])
    defparam i1_4_lut_adj_341.init = 16'hefff;
    LUT4 n946_bdd_2_lut_35027_rep_1049_3_lut (.A(n42801), .B(n45105), .C(n41229), 
         .Z(n45069)) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam n946_bdd_2_lut_35027_rep_1049_3_lut.init = 16'hb0b0;
    LUT4 i1_4_lut_adj_342 (.A(n34912), .B(n30136), .C(x_result_sel_csr_d), 
         .D(n34570), .Z(n34578)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(402[14:76])
    defparam i1_4_lut_adj_342.init = 16'hfff7;
    LUT4 i1_4_lut_adj_343 (.A(n31427), .B(n41213), .C(n41214), .D(n6781), 
         .Z(n34570)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(402[14:76])
    defparam i1_4_lut_adj_343.init = 16'hffdf;
    LUT4 i1_2_lut_rep_1003 (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .Z(n41408)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut_rep_1003.init = 16'hdddd;
    LUT4 i1_2_lut_3_lut (.A(\genblk1.wait_one_tick_done ), .B(n6781), .C(n6760), 
         .Z(n2)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_4_lut_adj_344 (.A(n34912), .B(n19987), .C(n30136), .D(n34908), 
         .Z(n31549)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_344.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_adj_345 (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n6761), .Z(n2_adj_146)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_345.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_346 (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n6762), .Z(n2_adj_147)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_346.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_347 (.A(\genblk1.wait_one_tick_done ), .B(n6781), 
         .C(n6763), .Z(n2_adj_148)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_347.init = 16'h2020;
    LUT4 i25263_4_lut (.A(n41241), .B(n41295), .C(n30216), .D(n31505), 
         .Z(m_result_sel_compare_d)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(402[14:76])
    defparam i25263_4_lut.init = 16'ha0a8;
    LUT4 i1_3_lut_4_lut_adj_348 (.A(n45105), .B(n41451), .C(n41452), .D(n41296), 
         .Z(n30058)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;
    defparam i1_3_lut_4_lut_adj_348.init = 16'hd000;
    LUT4 i1_4_lut_adj_349 (.A(n6775), .B(n6780), .C(n6777), .D(n6776), 
         .Z(n31829)) /* synthesis lut_function=(!(A+(B+!(C (D)+!C !(D))))) */ ;
    defparam i1_4_lut_adj_349.init = 16'h1001;
    LUT4 i5247_3_lut_4_lut (.A(n6780), .B(n41382), .C(n6768), .D(n6764), 
         .Z(n10589)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i5247_3_lut_4_lut.init = 16'hf780;
    LUT4 n40093_bdd_3_lut_4_lut (.A(n6780), .B(n41382), .C(n45183), .D(n40093), 
         .Z(n40094)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n40093_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i5243_3_lut_4_lut (.A(n6780), .B(n41382), .C(n6766), .D(n6764), 
         .Z(n10585)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i5243_3_lut_4_lut.init = 16'hf780;
    LUT4 i5249_3_lut_4_lut (.A(n6780), .B(n41382), .C(n6769), .D(n6764), 
         .Z(n10591)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i5249_3_lut_4_lut.init = 16'hf780;
    LUT4 i5139_2_lut_rep_1014 (.A(n6778), .B(n6779), .Z(n41419)) /* synthesis lut_function=(A+(B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(374[20:65])
    defparam i5139_2_lut_rep_1014.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut_adj_350 (.A(n6778), .B(n6779), .C(n6781), 
         .D(\genblk1.wait_one_tick_done ), .Z(n33940)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(374[20:65])
    defparam i1_2_lut_3_lut_4_lut_adj_350.init = 16'h0e00;
    LUT4 i5143_2_lut_3_lut_4_lut (.A(n6778), .B(n6779), .C(n10475), .D(n6777), 
         .Z(n10485)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(374[20:65])
    defparam i5143_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i5141_2_lut_rep_914_3_lut (.A(n6778), .B(n6779), .C(n6777), .Z(n41319)) /* synthesis lut_function=(A+(B+(C))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(374[20:65])
    defparam i5141_2_lut_rep_914_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_351 (.A(n41227), .B(n41363), .C(x_bypass_enable_x), 
         .D(n31542), .Z(n32006)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A (C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_351.init = 16'h080f;
    LUT4 i1_2_lut_3_lut_4_lut_adj_352 (.A(n41227), .B(n41363), .C(m_bypass_enable_m), 
         .D(n31542), .Z(n31984)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A (C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_352.init = 16'h080f;
    LUT4 i5251_3_lut_4_lut (.A(n6780), .B(n41382), .C(n6770), .D(n6764), 
         .Z(n10593)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i5251_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_3_lut_4_lut_adj_353 (.A(n41287), .B(n41229), .C(n41280), .D(n30820), 
         .Z(n35016)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(395[20:70])
    defparam i1_3_lut_4_lut_adj_353.init = 16'he000;
    LUT4 i5245_3_lut_4_lut (.A(n6780), .B(n41382), .C(n6767), .D(n6764), 
         .Z(n10587)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i5245_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_1033 (.A(n6780), .B(n6781), .Z(n41438)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut_rep_1033.init = 16'hdddd;
    LUT4 i1_2_lut_rep_907_3_lut (.A(n6780), .B(n6781), .C(n45105), .Z(n41312)) /* synthesis lut_function=((B+!(C))+!A) */ ;
    defparam i1_2_lut_rep_907_3_lut.init = 16'hdfdf;
    LUT4 i1_3_lut_4_lut_4_lut_adj_354 (.A(n6780), .B(n6781), .C(n41439), 
         .D(n41437), .Z(n35086)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_354.init = 16'hfffd;
    LUT4 i1_3_lut_rep_1034 (.A(\genblk1.wait_one_tick_done ), .B(n6778), 
         .C(n6781), .Z(n41439)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_rep_1034.init = 16'hf7f7;
    LUT4 i1_4_lut_4_lut (.A(\genblk1.wait_one_tick_done ), .B(n6778), .C(n6781), 
         .D(n10479), .Z(n35068)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_4_lut_4_lut.init = 16'hfff7;
    LUT4 i1_2_lut_rep_1035 (.A(n6779), .B(n6781), .Z(n41440)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut_rep_1035.init = 16'hdddd;
    LUT4 i1_3_lut_rep_959_4_lut (.A(n6779), .B(n6781), .C(n6780), .D(\genblk1.wait_one_tick_done ), 
         .Z(n41364)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;
    defparam i1_3_lut_rep_959_4_lut.init = 16'hdfff;
    LUT4 i1_2_lut_3_lut_adj_355 (.A(n6779), .B(n6781), .C(n45106), .Z(n32356)) /* synthesis lut_function=((B+!(C))+!A) */ ;
    defparam i1_2_lut_3_lut_adj_355.init = 16'hdfdf;
    LUT4 i1_3_lut_rep_1036 (.A(n45105), .B(n6777), .C(n6781), .Z(n41441)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_rep_1036.init = 16'hf7f7;
    LUT4 i1_2_lut_rep_881_3_lut_4_lut_4_lut (.A(\genblk1.wait_one_tick_done ), 
         .B(n6777), .C(n6781), .D(n6775), .Z(n41286)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_rep_881_3_lut_4_lut_4_lut.init = 16'hfff7;
    LUT4 i1_3_lut_4_lut_adj_356 (.A(n41363), .B(n31542), .C(n41296), .D(n30820), 
         .Z(n34474)) /* synthesis lut_function=(A (C+!(D))+!A (B+(C+!(D)))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(347[20:68])
    defparam i1_3_lut_4_lut_adj_356.init = 16'hf4ff;
    LUT4 i33188_2_lut_rep_779_3_lut_4_lut (.A(n41363), .B(n31542), .C(n45069), 
         .D(n41281), .Z(n41184)) /* synthesis lut_function=(!(A (C+(D))+!A !(B+!(C+(D))))) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(347[20:68])
    defparam i33188_2_lut_rep_779_3_lut_4_lut.init = 16'h444f;
    LUT4 i1_rep_787_4_lut (.A(n41365), .B(n41296), .C(n32356), .D(n45069), 
         .Z(n41192)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_rep_787_4_lut.init = 16'hfffe;
    LUT4 i33134_rep_175_2_lut_3_lut_4_lut (.A(n34474), .B(n41208), .C(n45069), 
         .D(n41281), .Z(n37939)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i33134_rep_175_2_lut_3_lut_4_lut.init = 16'h4440;
    LUT4 i1_2_lut_rep_1046 (.A(n6775), .B(n6781), .Z(n41451)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut_rep_1046.init = 16'hdddd;
    LUT4 i1_2_lut_rep_889_3_lut (.A(n6775), .B(n6781), .C(\genblk1.wait_one_tick_done ), 
         .Z(n41294)) /* synthesis lut_function=((B+!(C))+!A) */ ;
    defparam i1_2_lut_rep_889_3_lut.init = 16'hdfdf;
    LUT4 i1_2_lut_3_lut_4_lut_adj_357 (.A(n41295), .B(n41367), .C(n35086), 
         .D(n41294), .Z(n11815)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(349[20:68])
    defparam i1_2_lut_3_lut_4_lut_adj_357.init = 16'hfffb;
    LUT4 i1_3_lut_4_lut_adj_358 (.A(n41295), .B(n41367), .C(n41366), .D(n41287), 
         .Z(n31675)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(349[20:68])
    defparam i1_3_lut_4_lut_adj_358.init = 16'hfffb;
    LUT4 i1_2_lut_rep_796_3_lut_4_lut (.A(n41295), .B(n41367), .C(n11807), 
         .D(n41294), .Z(n41201)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(349[20:68])
    defparam i1_2_lut_rep_796_3_lut_4_lut.init = 16'hfffb;
    LUT4 i1_4_lut_4_lut_4_lut (.A(n6775), .B(n6781), .C(n10487), .D(n45106), 
         .Z(n11834)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam i1_4_lut_4_lut_4_lut.init = 16'hfdff;
    LUT4 instruction_30__I_0_172_i6_2_lut_rep_839_3_lut_3_lut_4_lut_4_lut (.A(n6775), 
         .B(n6781), .C(\genblk1.wait_one_tick_done ), .D(n6776), .Z(n41244)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam instruction_30__I_0_172_i6_2_lut_rep_839_3_lut_3_lut_4_lut_4_lut.init = 16'hffdf;
    LUT4 i15182_2_lut_rep_799_3_lut_4_lut (.A(n41441), .B(n41366), .C(n41363), 
         .D(n41367), .Z(n41204)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;
    defparam i15182_2_lut_rep_799_3_lut_4_lut.init = 16'he0f0;
    LUT4 i33134_2_lut_3_lut_4_lut (.A(n34474), .B(n41208), .C(n45069), 
         .D(n41281), .Z(\d_result_sel_1_d[1] )) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i33134_2_lut_3_lut_4_lut.init = 16'h4440;
    LUT4 i5253_3_lut_4_lut (.A(n6780), .B(n41382), .C(n6771), .D(n6764), 
         .Z(n10595)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i5253_3_lut_4_lut.init = 16'hf780;
    LUT4 i33134_rep_169_2_lut_3_lut_4_lut (.A(n34474), .B(n41208), .C(n45069), 
         .D(n41281), .Z(n37933)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i33134_rep_169_2_lut_3_lut_4_lut.init = 16'h4440;
    LUT4 i33160_2_lut_rep_800_3_lut_4_lut (.A(n41441), .B(n41366), .C(n41287), 
         .D(n41367), .Z(n41205)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i33160_2_lut_rep_800_3_lut_4_lut.init = 16'h0001;
    LUT4 i33110_2_lut_3_lut_4_lut (.A(n41441), .B(n41366), .C(n11807), 
         .D(n41367), .Z(x_result_sel_csr_d)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i33110_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i33134_rep_170_2_lut_3_lut_4_lut (.A(n34474), .B(n41208), .C(n45069), 
         .D(n41281), .Z(n37934)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i33134_rep_170_2_lut_3_lut_4_lut.init = 16'h4440;
    LUT4 i33134_rep_172_2_lut_3_lut_4_lut (.A(n34474), .B(n41208), .C(n45069), 
         .D(n41281), .Z(n37936)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i33134_rep_172_2_lut_3_lut_4_lut.init = 16'h4440;
    LUT4 i5115_3_lut_4_lut (.A(n6780), .B(n41382), .C(n6765), .D(n6764), 
         .Z(n10452)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i5115_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_rep_886 (.A(n41408), .B(n41365), .C(n41362), .D(n31829), 
         .Z(n41291)) /* synthesis lut_function=(A (B (C))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_rep_886.init = 16'hc080;
    LUT4 i33134_rep_173_2_lut_3_lut_4_lut (.A(n34474), .B(n41208), .C(n45069), 
         .D(n41281), .Z(n37937)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i33134_rep_173_2_lut_3_lut_4_lut.init = 16'h4440;
    LUT4 i33134_rep_174_2_lut_3_lut_4_lut (.A(n34474), .B(n41208), .C(n45069), 
         .D(n41281), .Z(n37938)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i33134_rep_174_2_lut_3_lut_4_lut.init = 16'h4440;
    LUT4 i33134_rep_171_2_lut_3_lut_4_lut (.A(n34474), .B(n41208), .C(n45069), 
         .D(n41281), .Z(n37935)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i33134_rep_171_2_lut_3_lut_4_lut.init = 16'h4440;
    LUT4 i2_4_lut_else_3_lut (.A(n45075), .B(\genblk1.wait_one_tick_done ), 
         .C(n6781), .D(n6776), .Z(n41462)) /* synthesis lut_function=(A+!((C+!(D))+!B)) */ ;
    defparam i2_4_lut_else_3_lut.init = 16'haeaa;
    LUT4 i1_3_lut_adj_359 (.A(n19987), .B(n19888), .C(n6028), .Z(n31494)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i1_3_lut_adj_359.init = 16'h0202;
    
endmodule
//
// Verilog Description of module lm32_adder
//

module lm32_adder (operand_0_x, operand_1_x, adder_op_x, adder_op_x_n, 
            adder_result_x, adder_carry_n_x) /* synthesis syn_module_defined=1 */ ;
    input [31:0]operand_0_x;
    input [31:0]operand_1_x;
    input adder_op_x;
    input adder_op_x_n;
    output [31:0]adder_result_x;
    output adder_carry_n_x;
    
    
    lm32_addsub addsub (.operand_0_x({operand_0_x}), .operand_1_x({operand_1_x}), 
            .adder_op_x(adder_op_x), .adder_op_x_n(adder_op_x_n), .adder_result_x({adder_result_x}), 
            .adder_carry_n_x(adder_carry_n_x)) /* synthesis syn_module_defined=1 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_adder.v(100[13] 109[6])
    
endmodule
//
// Verilog Description of module lm32_addsub
//

module lm32_addsub (operand_0_x, operand_1_x, adder_op_x, adder_op_x_n, 
            adder_result_x, adder_carry_n_x) /* synthesis syn_module_defined=1 */ ;
    input [31:0]operand_0_x;
    input [31:0]operand_1_x;
    input adder_op_x;
    input adder_op_x_n;
    output [31:0]adder_result_x;
    output adder_carry_n_x;
    
    
    pmi_addsubEo3232491b9e8 pmi_addsubECP5Uoff3232 (.DataA({operand_0_x}), 
            .DataB({operand_1_x}), .Result({adder_result_x}), .Cin(adder_op_x), 
            .Add_Sub(adder_op_x_n), .Cout(adder_carry_n_x)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=16, LSE_LCOL=13, LSE_RCOL=6, LSE_LLINE=100, LSE_RLINE=109 */ ;   // D:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/lm32_top/rtl/verilog/lm32_adder.v(100[13] 109[6])
    defparam pmi_addsubECP5Uoff3232.module_type = "pmi_addsub";
    defparam pmi_addsubECP5Uoff3232.pmi_family = "ECP5U";
    defparam pmi_addsubECP5Uoff3232.pmi_sign = "off";
    defparam pmi_addsubECP5Uoff3232.pmi_result_width = 32;
    defparam pmi_addsubECP5Uoff3232.pmi_data_width = 32;
    
endmodule
//
// Verilog Description of module \gpio(DATA_WIDTH=32'b01000,INPUT_WIDTH=32'b01,OUTPUT_WIDTH=32'b01,EDGE=1,POSE_EDGE_IRQ=1,INPUT_PORTS_ONLY=0,OUTPUT_PORTS_ONLY=1) 
//

module \gpio(DATA_WIDTH=32'b01000,INPUT_WIDTH=32'b01,OUTPUT_WIDTH=32'b01,EDGE=1,POSE_EDGE_IRQ=1,INPUT_PORTS_ONLY=0,OUTPUT_PORTS_ONLY=1)  (LEDGPIO_ACK_O, 
            REF_CLK_c, REF_CLK_c_enable_1606, PIO_OUT_7__N_3493, LED_R_c_0, 
            REF_CLK_c_enable_424, n36338, n41345, n41344, write_ack_N_4033, 
            n41185, n30156, n41347, dw10_cs_N_4471, dw00_cs_N_4467) /* synthesis syn_module_defined=1 */ ;
    output LEDGPIO_ACK_O;
    input REF_CLK_c;
    input REF_CLK_c_enable_1606;
    input PIO_OUT_7__N_3493;
    output LED_R_c_0;
    input REF_CLK_c_enable_424;
    input n36338;
    input n41345;
    input n41344;
    input write_ack_N_4033;
    output n41185;
    input n30156;
    input n41347;
    output dw10_cs_N_4471;
    output dw00_cs_N_4467;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    
    FD1S3DX GPIO_ACK_O_181 (.D(PIO_OUT_7__N_3493), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(LEDGPIO_ACK_O)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=638, LSE_RLINE=654 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/gpio/rtl/verilog/gpio.v(188[11] 191[33])
    defparam GPIO_ACK_O_181.GSR = "ENABLED";
    FD1P3DX PIO_DATA_0__182 (.D(n36338), .SP(REF_CLK_c_enable_424), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(LED_R_c_0)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=638, LSE_RLINE=654 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/gpio/rtl/verilog/gpio.v(258[11] 259[62])
    defparam PIO_DATA_0__182.GSR = "ENABLED";
    LUT4 write_ack_N_4033_I_0_132_2_lut_rep_780_3_lut (.A(n41345), .B(n41344), 
         .C(write_ack_N_4033), .Z(n41185)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/gpio/rtl/verilog/gpio.v(180[20:44])
    defparam write_ack_N_4033_I_0_132_2_lut_rep_780_3_lut.init = 16'h1010;
    LUT4 i33331_3_lut_4_lut (.A(n41345), .B(n41344), .C(n30156), .D(n41347), 
         .Z(dw10_cs_N_4471)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/gpio/rtl/verilog/gpio.v(180[20:44])
    defparam i33331_3_lut_4_lut.init = 16'h0100;
    LUT4 i33116_2_lut_3_lut_4_lut (.A(n41345), .B(n41344), .C(n30156), 
         .D(n41347), .Z(dw00_cs_N_4467)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/gpio/rtl/verilog/gpio.v(180[20:44])
    defparam i33116_2_lut_3_lut_4_lut.init = 16'h0001;
    
endmodule
//
// Verilog Description of module \Reg_Comp(reg_08_int_val=32'b010010001101001010101111001101,CLK_MHZ=48.0) 
//

module \Reg_Comp(reg_08_int_val=32'b010010001101001010101111001101,CLK_MHZ=48.0)  (LED_G_c_0, 
            REF_CLK_c, REF_CLK_c_enable_1606, n41328, \reg_04[0] , write_ack, 
            n35736, n15, n41301, n31750, n41210, n41303, n35854, 
            n41273, n41260, n35739, n41235, \SHAREDBUS_ADR_I[22] , 
            \SHAREDBUS_ADR_I[29] , write_ack_N_4033, n41251, n41324, 
            n41243, n41238, n41309, n41239, n41329, \GPOout_pins[2] , 
            n41330, \GPOout_pins[3] , n41331, \GPOout_pins[4] , n41332, 
            n41333, \GPOout_pins[6] , n41334, \GPOout_pins[7] , n41335, 
            \SHAREDBUS_DAT_I[8] , \reg_00[9] , \SHAREDBUS_DAT_I[9] , \SHAREDBUS_DAT_I[10] , 
            \reg_00[11] , \SHAREDBUS_DAT_I[11] , \SHAREDBUS_DAT_I[12] , 
            \reg_00[13] , \SHAREDBUS_DAT_I[13] , \reg_00[14] , \SHAREDBUS_DAT_I[14] , 
            \reg_00[15] , \SHAREDBUS_DAT_I[15] , n41336, \reg_00[17] , 
            n41337, \reg_00[18] , n41338, n41339, n41340, \reg_00[21] , 
            n41341, \reg_00[22] , n41342, n41343, \reg_00[24] , \SHAREDBUS_DAT_I[24] , 
            \reg_00[25] , \SHAREDBUS_DAT_I[25] , \SHAREDBUS_DAT_I[26] , 
            \SHAREDBUS_DAT_I[27] , \reg_00[28] , \SHAREDBUS_DAT_I[28] , 
            \reg_00[29] , \SHAREDBUS_DAT_I[29] , \SHAREDBUS_DAT_I[30] , 
            \SHAREDBUS_DAT_I[31] , n41279, n13, n13_adj_138, n13_adj_139, 
            n9, \reg_04[2] , \reg_04[3] , \reg_04[4] , \reg_04[6] , 
            \reg_04[7] , \reg_04[9] , \reg_04[11] , \reg_04[13] , \reg_04[14] , 
            \reg_04[15] , \reg_04[17] , \reg_04[18] , \reg_04[21] , 
            \reg_04[22] , \reg_04[24] , \reg_04[25] , \reg_04[28] , 
            \reg_04[29] , \GPOwb_DAT_O[8] , \GPOwb_DAT_O[1] , n13_adj_140, 
            n13_adj_141, n34304, n41185, n34112, \GPOwb_DAT_O[0] , 
            n11, n13_adj_142, \GPOwb_DAT_O[5] , n13_adj_143, n13_adj_144, 
            \SHAREDBUS_ADR_I[20] , n41242, n41250, n35577, n32366, 
            n41310, n19, n41225, n35647, n41258, n35724, n41253, 
            n41246, \SHAREDBUS_ADR_I[26] , \SHAREDBUS_ADR_I[16] , n35633, 
            read_ack, n41269, n34242, n41304, n33328, n33294, n32312, 
            n33404, n33370, n33290, \SHAREDBUS_ADR_I[24] , \SHAREDBUS_ADR_I[25] , 
            \SHAREDBUS_ADR_I[18] , \SHAREDBUS_ADR_I[27] , n33256, n33252, 
            n33218, n33214, n33180, n33356, n33366) /* synthesis syn_module_defined=1 */ ;
    output LED_G_c_0;
    input REF_CLK_c;
    input REF_CLK_c_enable_1606;
    input n41328;
    output \reg_04[0] ;
    output write_ack;
    input n35736;
    input n15;
    input n41301;
    output n31750;
    input n41210;
    input n41303;
    input n35854;
    output n41273;
    output n41260;
    output n35739;
    input n41235;
    input \SHAREDBUS_ADR_I[22] ;
    input \SHAREDBUS_ADR_I[29] ;
    output write_ack_N_4033;
    input n41251;
    input n41324;
    input n41243;
    input n41238;
    input n41309;
    input n41239;
    input n41329;
    output \GPOout_pins[2] ;
    input n41330;
    output \GPOout_pins[3] ;
    input n41331;
    output \GPOout_pins[4] ;
    input n41332;
    input n41333;
    output \GPOout_pins[6] ;
    input n41334;
    output \GPOout_pins[7] ;
    input n41335;
    input \SHAREDBUS_DAT_I[8] ;
    output \reg_00[9] ;
    input \SHAREDBUS_DAT_I[9] ;
    input \SHAREDBUS_DAT_I[10] ;
    output \reg_00[11] ;
    input \SHAREDBUS_DAT_I[11] ;
    input \SHAREDBUS_DAT_I[12] ;
    output \reg_00[13] ;
    input \SHAREDBUS_DAT_I[13] ;
    output \reg_00[14] ;
    input \SHAREDBUS_DAT_I[14] ;
    output \reg_00[15] ;
    input \SHAREDBUS_DAT_I[15] ;
    input n41336;
    output \reg_00[17] ;
    input n41337;
    output \reg_00[18] ;
    input n41338;
    input n41339;
    input n41340;
    output \reg_00[21] ;
    input n41341;
    output \reg_00[22] ;
    input n41342;
    input n41343;
    output \reg_00[24] ;
    input \SHAREDBUS_DAT_I[24] ;
    output \reg_00[25] ;
    input \SHAREDBUS_DAT_I[25] ;
    input \SHAREDBUS_DAT_I[26] ;
    input \SHAREDBUS_DAT_I[27] ;
    output \reg_00[28] ;
    input \SHAREDBUS_DAT_I[28] ;
    output \reg_00[29] ;
    input \SHAREDBUS_DAT_I[29] ;
    input \SHAREDBUS_DAT_I[30] ;
    input \SHAREDBUS_DAT_I[31] ;
    input n41279;
    output n13;
    output n13_adj_138;
    output n13_adj_139;
    output n9;
    output \reg_04[2] ;
    output \reg_04[3] ;
    output \reg_04[4] ;
    output \reg_04[6] ;
    output \reg_04[7] ;
    output \reg_04[9] ;
    output \reg_04[11] ;
    output \reg_04[13] ;
    output \reg_04[14] ;
    output \reg_04[15] ;
    output \reg_04[17] ;
    output \reg_04[18] ;
    output \reg_04[21] ;
    output \reg_04[22] ;
    output \reg_04[24] ;
    output \reg_04[25] ;
    output \reg_04[28] ;
    output \reg_04[29] ;
    output \GPOwb_DAT_O[8] ;
    output \GPOwb_DAT_O[1] ;
    output n13_adj_140;
    output n13_adj_141;
    input n34304;
    input n41185;
    input n34112;
    output \GPOwb_DAT_O[0] ;
    output n11;
    output n13_adj_142;
    output \GPOwb_DAT_O[5] ;
    output n13_adj_143;
    output n13_adj_144;
    input \SHAREDBUS_ADR_I[20] ;
    output n41242;
    input n41250;
    input n35577;
    input n32366;
    input n41310;
    input n19;
    input n41225;
    input n35647;
    input n41258;
    input n35724;
    input n41253;
    input n41246;
    input \SHAREDBUS_ADR_I[26] ;
    input \SHAREDBUS_ADR_I[16] ;
    input n35633;
    output read_ack;
    input n41269;
    input n34242;
    input n41304;
    output n33328;
    input n33294;
    input n32312;
    output n33404;
    input n33370;
    output n33290;
    input \SHAREDBUS_ADR_I[24] ;
    input \SHAREDBUS_ADR_I[25] ;
    input \SHAREDBUS_ADR_I[18] ;
    input \SHAREDBUS_ADR_I[27] ;
    input n33256;
    output n33252;
    input n33218;
    output n33214;
    input n33180;
    input n33356;
    output n33366;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    
    \wb_reg_dev(CLK_MHZ=48.0)  instantiate_wb_reg_dev (.LED_G_c_0(LED_G_c_0), 
            .REF_CLK_c(REF_CLK_c), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .n41328(n41328), .reg_04({Open_73, Open_74, Open_75, Open_76, 
            Open_77, Open_78, Open_79, Open_80, Open_81, Open_82, 
            Open_83, Open_84, Open_85, Open_86, Open_87, Open_88, 
            Open_89, Open_90, Open_91, Open_92, Open_93, Open_94, 
            Open_95, Open_96, Open_97, Open_98, Open_99, Open_100, 
            Open_101, Open_102, Open_103, \reg_04[0] }), .write_ack(write_ack), 
            .n35736(n35736), .n15(n15), .n41301(n41301), .n31750(n31750), 
            .n41210(n41210), .n41303(n41303), .n35854(n35854), .n41273(n41273), 
            .n41260(n41260), .n35739(n35739), .n41235(n41235), .\SHAREDBUS_ADR_I[22] (\SHAREDBUS_ADR_I[22] ), 
            .\SHAREDBUS_ADR_I[29] (\SHAREDBUS_ADR_I[29] ), .write_ack_N_4033(write_ack_N_4033), 
            .n41251(n41251), .n41324(n41324), .n41243(n41243), .n41238(n41238), 
            .n41309(n41309), .n41239(n41239), .n41329(n41329), .\GPOout_pins[2] (\GPOout_pins[2] ), 
            .n41330(n41330), .\GPOout_pins[3] (\GPOout_pins[3] ), .n41331(n41331), 
            .\GPOout_pins[4] (\GPOout_pins[4] ), .n41332(n41332), .n41333(n41333), 
            .\GPOout_pins[6] (\GPOout_pins[6] ), .n41334(n41334), .\GPOout_pins[7] (\GPOout_pins[7] ), 
            .n41335(n41335), .\SHAREDBUS_DAT_I[8] (\SHAREDBUS_DAT_I[8] ), 
            .\reg_00[9] (\reg_00[9] ), .\SHAREDBUS_DAT_I[9] (\SHAREDBUS_DAT_I[9] ), 
            .\SHAREDBUS_DAT_I[10] (\SHAREDBUS_DAT_I[10] ), .\reg_00[11] (\reg_00[11] ), 
            .\SHAREDBUS_DAT_I[11] (\SHAREDBUS_DAT_I[11] ), .\SHAREDBUS_DAT_I[12] (\SHAREDBUS_DAT_I[12] ), 
            .\reg_00[13] (\reg_00[13] ), .\SHAREDBUS_DAT_I[13] (\SHAREDBUS_DAT_I[13] ), 
            .\reg_00[14] (\reg_00[14] ), .\SHAREDBUS_DAT_I[14] (\SHAREDBUS_DAT_I[14] ), 
            .\reg_00[15] (\reg_00[15] ), .\SHAREDBUS_DAT_I[15] (\SHAREDBUS_DAT_I[15] ), 
            .n41336(n41336), .\reg_00[17] (\reg_00[17] ), .n41337(n41337), 
            .\reg_00[18] (\reg_00[18] ), .n41338(n41338), .n41339(n41339), 
            .n41340(n41340), .\reg_00[21] (\reg_00[21] ), .n41341(n41341), 
            .\reg_00[22] (\reg_00[22] ), .n41342(n41342), .n41343(n41343), 
            .\reg_00[24] (\reg_00[24] ), .\SHAREDBUS_DAT_I[24] (\SHAREDBUS_DAT_I[24] ), 
            .\reg_00[25] (\reg_00[25] ), .\SHAREDBUS_DAT_I[25] (\SHAREDBUS_DAT_I[25] ), 
            .\SHAREDBUS_DAT_I[26] (\SHAREDBUS_DAT_I[26] ), .\SHAREDBUS_DAT_I[27] (\SHAREDBUS_DAT_I[27] ), 
            .\reg_00[28] (\reg_00[28] ), .\SHAREDBUS_DAT_I[28] (\SHAREDBUS_DAT_I[28] ), 
            .\reg_00[29] (\reg_00[29] ), .\SHAREDBUS_DAT_I[29] (\SHAREDBUS_DAT_I[29] ), 
            .\SHAREDBUS_DAT_I[30] (\SHAREDBUS_DAT_I[30] ), .\SHAREDBUS_DAT_I[31] (\SHAREDBUS_DAT_I[31] ), 
            .n41279(n41279), .n13(n13), .n13_adj_131(n13_adj_138), .n13_adj_132(n13_adj_139), 
            .n9(n9), .\reg_04[2] (\reg_04[2] ), .\reg_04[3] (\reg_04[3] ), 
            .\reg_04[4] (\reg_04[4] ), .\reg_04[6] (\reg_04[6] ), .\reg_04[7] (\reg_04[7] ), 
            .\reg_04[9] (\reg_04[9] ), .\reg_04[11] (\reg_04[11] ), .\reg_04[13] (\reg_04[13] ), 
            .\reg_04[14] (\reg_04[14] ), .\reg_04[15] (\reg_04[15] ), .\reg_04[17] (\reg_04[17] ), 
            .\reg_04[18] (\reg_04[18] ), .\reg_04[21] (\reg_04[21] ), .\reg_04[22] (\reg_04[22] ), 
            .\reg_04[24] (\reg_04[24] ), .\reg_04[25] (\reg_04[25] ), .\reg_04[28] (\reg_04[28] ), 
            .\reg_04[29] (\reg_04[29] ), .\GPOwb_DAT_O[8] (\GPOwb_DAT_O[8] ), 
            .\GPOwb_DAT_O[1] (\GPOwb_DAT_O[1] ), .n13_adj_133(n13_adj_140), 
            .n13_adj_134(n13_adj_141), .n34304(n34304), .n41185(n41185), 
            .n34112(n34112), .\GPOwb_DAT_O[0] (\GPOwb_DAT_O[0] ), .n11(n11), 
            .n13_adj_135(n13_adj_142), .\GPOwb_DAT_O[5] (\GPOwb_DAT_O[5] ), 
            .n13_adj_136(n13_adj_143), .n13_adj_137(n13_adj_144), .\SHAREDBUS_ADR_I[20] (\SHAREDBUS_ADR_I[20] ), 
            .n41242(n41242), .n41250(n41250), .n35577(n35577), .n32366(n32366), 
            .n41310(n41310), .n19(n19), .n41225(n41225), .n35647(n35647), 
            .n41258(n41258), .n35724(n35724), .n41253(n41253), .n41246(n41246), 
            .\SHAREDBUS_ADR_I[26] (\SHAREDBUS_ADR_I[26] ), .\SHAREDBUS_ADR_I[16] (\SHAREDBUS_ADR_I[16] ), 
            .n35633(n35633), .read_ack(read_ack), .n41269(n41269), .n34242(n34242), 
            .n41304(n41304), .n33328(n33328), .n33294(n33294), .n32312(n32312), 
            .n33404(n33404), .n33370(n33370), .n33290(n33290), .\SHAREDBUS_ADR_I[24] (\SHAREDBUS_ADR_I[24] ), 
            .\SHAREDBUS_ADR_I[25] (\SHAREDBUS_ADR_I[25] ), .\SHAREDBUS_ADR_I[18] (\SHAREDBUS_ADR_I[18] ), 
            .\SHAREDBUS_ADR_I[27] (\SHAREDBUS_ADR_I[27] ), .n33256(n33256), 
            .n33252(n33252), .n33218(n33218), .n33214(n33214), .n33180(n33180), 
            .n33356(n33356), .n33366(n33366)) /* synthesis syn_module_defined=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/Reg_Comp.v(78[11] 97[34])
    
endmodule
//
// Verilog Description of module \wb_reg_dev(CLK_MHZ=48.0) 
//

module \wb_reg_dev(CLK_MHZ=48.0)  (LED_G_c_0, REF_CLK_c, REF_CLK_c_enable_1606, 
            n41328, reg_04, write_ack, n35736, n15, n41301, n31750, 
            n41210, n41303, n35854, n41273, n41260, n35739, n41235, 
            \SHAREDBUS_ADR_I[22] , \SHAREDBUS_ADR_I[29] , write_ack_N_4033, 
            n41251, n41324, n41243, n41238, n41309, n41239, n41329, 
            \GPOout_pins[2] , n41330, \GPOout_pins[3] , n41331, \GPOout_pins[4] , 
            n41332, n41333, \GPOout_pins[6] , n41334, \GPOout_pins[7] , 
            n41335, \SHAREDBUS_DAT_I[8] , \reg_00[9] , \SHAREDBUS_DAT_I[9] , 
            \SHAREDBUS_DAT_I[10] , \reg_00[11] , \SHAREDBUS_DAT_I[11] , 
            \SHAREDBUS_DAT_I[12] , \reg_00[13] , \SHAREDBUS_DAT_I[13] , 
            \reg_00[14] , \SHAREDBUS_DAT_I[14] , \reg_00[15] , \SHAREDBUS_DAT_I[15] , 
            n41336, \reg_00[17] , n41337, \reg_00[18] , n41338, n41339, 
            n41340, \reg_00[21] , n41341, \reg_00[22] , n41342, n41343, 
            \reg_00[24] , \SHAREDBUS_DAT_I[24] , \reg_00[25] , \SHAREDBUS_DAT_I[25] , 
            \SHAREDBUS_DAT_I[26] , \SHAREDBUS_DAT_I[27] , \reg_00[28] , 
            \SHAREDBUS_DAT_I[28] , \reg_00[29] , \SHAREDBUS_DAT_I[29] , 
            \SHAREDBUS_DAT_I[30] , \SHAREDBUS_DAT_I[31] , n41279, n13, 
            n13_adj_131, n13_adj_132, n9, \reg_04[2] , \reg_04[3] , 
            \reg_04[4] , \reg_04[6] , \reg_04[7] , \reg_04[9] , \reg_04[11] , 
            \reg_04[13] , \reg_04[14] , \reg_04[15] , \reg_04[17] , 
            \reg_04[18] , \reg_04[21] , \reg_04[22] , \reg_04[24] , 
            \reg_04[25] , \reg_04[28] , \reg_04[29] , \GPOwb_DAT_O[8] , 
            \GPOwb_DAT_O[1] , n13_adj_133, n13_adj_134, n34304, n41185, 
            n34112, \GPOwb_DAT_O[0] , n11, n13_adj_135, \GPOwb_DAT_O[5] , 
            n13_adj_136, n13_adj_137, \SHAREDBUS_ADR_I[20] , n41242, 
            n41250, n35577, n32366, n41310, n19, n41225, n35647, 
            n41258, n35724, n41253, n41246, \SHAREDBUS_ADR_I[26] , 
            \SHAREDBUS_ADR_I[16] , n35633, read_ack, n41269, n34242, 
            n41304, n33328, n33294, n32312, n33404, n33370, n33290, 
            \SHAREDBUS_ADR_I[24] , \SHAREDBUS_ADR_I[25] , \SHAREDBUS_ADR_I[18] , 
            \SHAREDBUS_ADR_I[27] , n33256, n33252, n33218, n33214, 
            n33180, n33356, n33366) /* synthesis syn_module_defined=1 */ ;
    output LED_G_c_0;
    input REF_CLK_c;
    input REF_CLK_c_enable_1606;
    input n41328;
    output [31:0]reg_04;
    output write_ack;
    input n35736;
    input n15;
    input n41301;
    output n31750;
    input n41210;
    input n41303;
    input n35854;
    output n41273;
    output n41260;
    output n35739;
    input n41235;
    input \SHAREDBUS_ADR_I[22] ;
    input \SHAREDBUS_ADR_I[29] ;
    output write_ack_N_4033;
    input n41251;
    input n41324;
    input n41243;
    input n41238;
    input n41309;
    input n41239;
    input n41329;
    output \GPOout_pins[2] ;
    input n41330;
    output \GPOout_pins[3] ;
    input n41331;
    output \GPOout_pins[4] ;
    input n41332;
    input n41333;
    output \GPOout_pins[6] ;
    input n41334;
    output \GPOout_pins[7] ;
    input n41335;
    input \SHAREDBUS_DAT_I[8] ;
    output \reg_00[9] ;
    input \SHAREDBUS_DAT_I[9] ;
    input \SHAREDBUS_DAT_I[10] ;
    output \reg_00[11] ;
    input \SHAREDBUS_DAT_I[11] ;
    input \SHAREDBUS_DAT_I[12] ;
    output \reg_00[13] ;
    input \SHAREDBUS_DAT_I[13] ;
    output \reg_00[14] ;
    input \SHAREDBUS_DAT_I[14] ;
    output \reg_00[15] ;
    input \SHAREDBUS_DAT_I[15] ;
    input n41336;
    output \reg_00[17] ;
    input n41337;
    output \reg_00[18] ;
    input n41338;
    input n41339;
    input n41340;
    output \reg_00[21] ;
    input n41341;
    output \reg_00[22] ;
    input n41342;
    input n41343;
    output \reg_00[24] ;
    input \SHAREDBUS_DAT_I[24] ;
    output \reg_00[25] ;
    input \SHAREDBUS_DAT_I[25] ;
    input \SHAREDBUS_DAT_I[26] ;
    input \SHAREDBUS_DAT_I[27] ;
    output \reg_00[28] ;
    input \SHAREDBUS_DAT_I[28] ;
    output \reg_00[29] ;
    input \SHAREDBUS_DAT_I[29] ;
    input \SHAREDBUS_DAT_I[30] ;
    input \SHAREDBUS_DAT_I[31] ;
    input n41279;
    output n13;
    output n13_adj_131;
    output n13_adj_132;
    output n9;
    output \reg_04[2] ;
    output \reg_04[3] ;
    output \reg_04[4] ;
    output \reg_04[6] ;
    output \reg_04[7] ;
    output \reg_04[9] ;
    output \reg_04[11] ;
    output \reg_04[13] ;
    output \reg_04[14] ;
    output \reg_04[15] ;
    output \reg_04[17] ;
    output \reg_04[18] ;
    output \reg_04[21] ;
    output \reg_04[22] ;
    output \reg_04[24] ;
    output \reg_04[25] ;
    output \reg_04[28] ;
    output \reg_04[29] ;
    output \GPOwb_DAT_O[8] ;
    output \GPOwb_DAT_O[1] ;
    output n13_adj_133;
    output n13_adj_134;
    input n34304;
    input n41185;
    input n34112;
    output \GPOwb_DAT_O[0] ;
    output n11;
    output n13_adj_135;
    output \GPOwb_DAT_O[5] ;
    output n13_adj_136;
    output n13_adj_137;
    input \SHAREDBUS_ADR_I[20] ;
    output n41242;
    input n41250;
    input n35577;
    input n32366;
    input n41310;
    input n19;
    input n41225;
    input n35647;
    input n41258;
    input n35724;
    input n41253;
    input n41246;
    input \SHAREDBUS_ADR_I[26] ;
    input \SHAREDBUS_ADR_I[16] ;
    input n35633;
    output read_ack;
    input n41269;
    input n34242;
    input n41304;
    output n33328;
    input n33294;
    input n32312;
    output n33404;
    input n33370;
    output n33290;
    input \SHAREDBUS_ADR_I[24] ;
    input \SHAREDBUS_ADR_I[25] ;
    input \SHAREDBUS_ADR_I[18] ;
    input \SHAREDBUS_ADR_I[27] ;
    input n33256;
    output n33252;
    input n33218;
    output n33214;
    input n33180;
    input n33356;
    output n33366;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    
    wire REF_CLK_c_enable_1487, REF_CLK_c_enable_1519, write_ack_N_4031, 
        n35944, n35926, REF_CLK_c_enable_1527, REF_CLK_c_enable_1535, 
        REF_CLK_c_enable_1543;
    wire [7:0]GPOout_pins;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1_vhd.vhd(11[3:14])
    wire [31:0]reg_00;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(80[15:21])
    
    wire REF_CLK_c_enable_1495, REF_CLK_c_enable_1503, REF_CLK_c_enable_1511;
    wire [31:0]reg_04_c;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(81[15:21])
    
    wire n18860, n18416, n18314, n18138;
    wire [31:0]wb_slave_data_31__N_3867;
    
    wire n18656, n18553, n18519, n18279, n18792, n18176, n32388, 
        n35914, n35820, n35128, n35894, n35112, n35583, n32110, 
        n35898, n32096, n33318, n35906, n35800, n33394, n33280, 
        n33242, n33204;
    
    FD1P3DX reg_00__i1 (.D(n41328), .SP(REF_CLK_c_enable_1487), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(LED_G_c_0)) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i1.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i0 (.D(n41328), .SP(REF_CLK_c_enable_1519), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_04[0])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i0.GSR = "ENABLED";
    FD1S3DX write_ack_125 (.D(write_ack_N_4031), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(write_ack)) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(125[12] 133[10])
    defparam write_ack_125.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n35736), .B(n15), .C(n35944), .D(n41301), .Z(n31750)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut.init = 16'h0100;
    LUT4 i30782_4_lut (.A(n41210), .B(n35926), .C(n41303), .D(n35854), 
         .Z(n35944)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i30782_4_lut.init = 16'hfffd;
    LUT4 i30764_4_lut (.A(n41273), .B(n41260), .C(n35739), .D(n41235), 
         .Z(n35926)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30764_4_lut.init = 16'hfffe;
    LUT4 i30579_2_lut (.A(\SHAREDBUS_ADR_I[22] ), .B(\SHAREDBUS_ADR_I[29] ), 
         .Z(n35739)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i30579_2_lut.init = 16'heeee;
    LUT4 i4226_2_lut_3_lut_4_lut (.A(write_ack_N_4033), .B(n41251), .C(n41324), 
         .D(n41243), .Z(REF_CLK_c_enable_1519)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(101[24] 102[31])
    defparam i4226_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i4919_2_lut_3_lut_4_lut (.A(write_ack_N_4033), .B(n41251), .C(n41238), 
         .D(n41243), .Z(REF_CLK_c_enable_1527)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(101[24] 102[31])
    defparam i4919_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i4935_2_lut_3_lut_4_lut (.A(write_ack_N_4033), .B(n41251), .C(n41309), 
         .D(n41243), .Z(REF_CLK_c_enable_1535)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(101[24] 102[31])
    defparam i4935_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i4951_2_lut_3_lut_4_lut (.A(write_ack_N_4033), .B(n41251), .C(n41239), 
         .D(n41243), .Z(REF_CLK_c_enable_1543)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(101[24] 102[31])
    defparam i4951_2_lut_3_lut_4_lut.init = 16'h2000;
    FD1P3DX reg_00__i2 (.D(n41329), .SP(REF_CLK_c_enable_1487), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(GPOout_pins[1])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i2.GSR = "ENABLED";
    FD1P3DX reg_00__i3 (.D(n41330), .SP(REF_CLK_c_enable_1487), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\GPOout_pins[2] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i3.GSR = "ENABLED";
    FD1P3DX reg_00__i4 (.D(n41331), .SP(REF_CLK_c_enable_1487), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\GPOout_pins[3] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i4.GSR = "ENABLED";
    FD1P3DX reg_00__i5 (.D(n41332), .SP(REF_CLK_c_enable_1487), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\GPOout_pins[4] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i5.GSR = "ENABLED";
    FD1P3DX reg_00__i6 (.D(n41333), .SP(REF_CLK_c_enable_1487), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(GPOout_pins[5])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i6.GSR = "ENABLED";
    FD1P3DX reg_00__i7 (.D(n41334), .SP(REF_CLK_c_enable_1487), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\GPOout_pins[6] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i7.GSR = "ENABLED";
    FD1P3DX reg_00__i8 (.D(n41335), .SP(REF_CLK_c_enable_1487), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\GPOout_pins[7] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i8.GSR = "ENABLED";
    FD1P3DX reg_00__i9 (.D(\SHAREDBUS_DAT_I[8] ), .SP(REF_CLK_c_enable_1495), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[8])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i9.GSR = "ENABLED";
    FD1P3DX reg_00__i10 (.D(\SHAREDBUS_DAT_I[9] ), .SP(REF_CLK_c_enable_1495), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_00[9] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i10.GSR = "ENABLED";
    FD1P3DX reg_00__i11 (.D(\SHAREDBUS_DAT_I[10] ), .SP(REF_CLK_c_enable_1495), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[10])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i11.GSR = "ENABLED";
    FD1P3DX reg_00__i12 (.D(\SHAREDBUS_DAT_I[11] ), .SP(REF_CLK_c_enable_1495), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_00[11] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i12.GSR = "ENABLED";
    FD1P3DX reg_00__i13 (.D(\SHAREDBUS_DAT_I[12] ), .SP(REF_CLK_c_enable_1495), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[12])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i13.GSR = "ENABLED";
    FD1P3DX reg_00__i14 (.D(\SHAREDBUS_DAT_I[13] ), .SP(REF_CLK_c_enable_1495), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_00[13] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i14.GSR = "ENABLED";
    FD1P3DX reg_00__i15 (.D(\SHAREDBUS_DAT_I[14] ), .SP(REF_CLK_c_enable_1495), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_00[14] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i15.GSR = "ENABLED";
    FD1P3DX reg_00__i16 (.D(\SHAREDBUS_DAT_I[15] ), .SP(REF_CLK_c_enable_1495), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_00[15] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i16.GSR = "ENABLED";
    FD1P3DX reg_00__i17 (.D(n41336), .SP(REF_CLK_c_enable_1503), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_00[16])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i17.GSR = "ENABLED";
    FD1P3DX reg_00__i18 (.D(n41337), .SP(REF_CLK_c_enable_1503), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_00[17] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i18.GSR = "ENABLED";
    FD1P3DX reg_00__i19 (.D(n41338), .SP(REF_CLK_c_enable_1503), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_00[18] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i19.GSR = "ENABLED";
    FD1P3DX reg_00__i20 (.D(n41339), .SP(REF_CLK_c_enable_1503), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_00[19])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i20.GSR = "ENABLED";
    FD1P3DX reg_00__i21 (.D(n41340), .SP(REF_CLK_c_enable_1503), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_00[20])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i21.GSR = "ENABLED";
    FD1P3DX reg_00__i22 (.D(n41341), .SP(REF_CLK_c_enable_1503), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_00[21] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i22.GSR = "ENABLED";
    FD1P3DX reg_00__i23 (.D(n41342), .SP(REF_CLK_c_enable_1503), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_00[22] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i23.GSR = "ENABLED";
    FD1P3DX reg_00__i24 (.D(n41343), .SP(REF_CLK_c_enable_1503), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_00[23])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i24.GSR = "ENABLED";
    FD1P3DX reg_00__i25 (.D(\SHAREDBUS_DAT_I[24] ), .SP(REF_CLK_c_enable_1511), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_00[24] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i25.GSR = "ENABLED";
    FD1P3DX reg_00__i26 (.D(\SHAREDBUS_DAT_I[25] ), .SP(REF_CLK_c_enable_1511), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_00[25] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i26.GSR = "ENABLED";
    FD1P3DX reg_00__i27 (.D(\SHAREDBUS_DAT_I[26] ), .SP(REF_CLK_c_enable_1511), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[26])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i27.GSR = "ENABLED";
    FD1P3DX reg_00__i28 (.D(\SHAREDBUS_DAT_I[27] ), .SP(REF_CLK_c_enable_1511), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[27])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i28.GSR = "ENABLED";
    FD1P3DX reg_00__i29 (.D(\SHAREDBUS_DAT_I[28] ), .SP(REF_CLK_c_enable_1511), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_00[28] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i29.GSR = "ENABLED";
    FD1P3DX reg_00__i30 (.D(\SHAREDBUS_DAT_I[29] ), .SP(REF_CLK_c_enable_1511), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_00[29] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i30.GSR = "ENABLED";
    FD1P3DX reg_00__i31 (.D(\SHAREDBUS_DAT_I[30] ), .SP(REF_CLK_c_enable_1511), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[30])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i31.GSR = "ENABLED";
    FD1P3DX reg_00__i32 (.D(\SHAREDBUS_DAT_I[31] ), .SP(REF_CLK_c_enable_1511), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[31])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(141[12] 157[10])
    defparam reg_00__i32.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i1 (.D(n41329), .SP(REF_CLK_c_enable_1519), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_04_c[1])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i1.GSR = "ENABLED";
    LUT4 i4997_2_lut_3_lut_4_lut (.A(write_ack_N_4033), .B(n41279), .C(n41309), 
         .D(n41243), .Z(REF_CLK_c_enable_1503)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(99[24] 100[31])
    defparam i4997_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i13578_3_lut_4_lut (.A(write_ack_N_4033), .B(n41279), .C(reg_00[10]), 
         .D(n18860), .Z(n13)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(99[24] 100[31])
    defparam i13578_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13121_3_lut_4_lut (.A(write_ack_N_4033), .B(n41279), .C(reg_00[23]), 
         .D(n18416), .Z(n13_adj_131)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(99[24] 100[31])
    defparam i13121_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13016_3_lut_4_lut (.A(write_ack_N_4033), .B(n41279), .C(reg_00[26]), 
         .D(n18314), .Z(n13_adj_132)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(99[24] 100[31])
    defparam i13016_3_lut_4_lut.init = 16'hfd20;
    LUT4 i12835_3_lut_4_lut (.A(write_ack_N_4033), .B(n41279), .C(reg_00[31]), 
         .D(n18138), .Z(n9)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(99[24] 100[31])
    defparam i12835_3_lut_4_lut.init = 16'hfd20;
    FD1P3DX reg_04_i0_i2 (.D(n41330), .SP(REF_CLK_c_enable_1519), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_04[2] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i2.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i3 (.D(n41331), .SP(REF_CLK_c_enable_1519), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_04[3] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i3.GSR = "ENABLED";
    FD1P3BX reg_04_i0_i4 (.D(n41332), .SP(REF_CLK_c_enable_1519), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(\reg_04[4] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i4.GSR = "ENABLED";
    FD1P3BX reg_04_i0_i5 (.D(n41333), .SP(REF_CLK_c_enable_1519), .CK(REF_CLK_c), 
            .PD(REF_CLK_c_enable_1606), .Q(reg_04_c[5])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i5.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i6 (.D(n41334), .SP(REF_CLK_c_enable_1519), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_04[6] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i6.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i7 (.D(n41335), .SP(REF_CLK_c_enable_1519), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_04[7] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i7.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i8 (.D(\SHAREDBUS_DAT_I[8] ), .SP(REF_CLK_c_enable_1527), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_04_c[8])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i8.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i9 (.D(\SHAREDBUS_DAT_I[9] ), .SP(REF_CLK_c_enable_1527), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_04[9] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i9.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i10 (.D(\SHAREDBUS_DAT_I[10] ), .SP(REF_CLK_c_enable_1527), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_04_c[10])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i10.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i11 (.D(\SHAREDBUS_DAT_I[11] ), .SP(REF_CLK_c_enable_1527), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_04[11] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i11.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i12 (.D(\SHAREDBUS_DAT_I[12] ), .SP(REF_CLK_c_enable_1527), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_04_c[12])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i12.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i13 (.D(\SHAREDBUS_DAT_I[13] ), .SP(REF_CLK_c_enable_1527), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_04[13] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i13.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i14 (.D(\SHAREDBUS_DAT_I[14] ), .SP(REF_CLK_c_enable_1527), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_04[14] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i14.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i15 (.D(\SHAREDBUS_DAT_I[15] ), .SP(REF_CLK_c_enable_1527), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_04[15] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i15.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i16 (.D(n41336), .SP(REF_CLK_c_enable_1535), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_04_c[16])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i16.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i17 (.D(n41337), .SP(REF_CLK_c_enable_1535), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_04[17] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i17.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i18 (.D(n41338), .SP(REF_CLK_c_enable_1535), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_04[18] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i18.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i19 (.D(n41339), .SP(REF_CLK_c_enable_1535), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_04_c[19])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i19.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i20 (.D(n41340), .SP(REF_CLK_c_enable_1535), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_04_c[20])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i20.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i21 (.D(n41341), .SP(REF_CLK_c_enable_1535), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_04[21] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i21.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i22 (.D(n41342), .SP(REF_CLK_c_enable_1535), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_04[22] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i22.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i23 (.D(n41343), .SP(REF_CLK_c_enable_1535), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_04_c[23])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i23.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i24 (.D(\SHAREDBUS_DAT_I[24] ), .SP(REF_CLK_c_enable_1543), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_04[24] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i24.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i25 (.D(\SHAREDBUS_DAT_I[25] ), .SP(REF_CLK_c_enable_1543), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_04[25] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i25.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i26 (.D(\SHAREDBUS_DAT_I[26] ), .SP(REF_CLK_c_enable_1543), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_04_c[26])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i26.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i27 (.D(\SHAREDBUS_DAT_I[27] ), .SP(REF_CLK_c_enable_1543), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_04_c[27])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i27.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i28 (.D(\SHAREDBUS_DAT_I[28] ), .SP(REF_CLK_c_enable_1543), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_04[28] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i28.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i29 (.D(\SHAREDBUS_DAT_I[29] ), .SP(REF_CLK_c_enable_1543), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_04[29] )) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i29.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i30 (.D(\SHAREDBUS_DAT_I[30] ), .SP(REF_CLK_c_enable_1543), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_04_c[30])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i30.GSR = "ENABLED";
    FD1P3DX reg_04_i0_i31 (.D(\SHAREDBUS_DAT_I[31] ), .SP(REF_CLK_c_enable_1543), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_04_c[31])) /* synthesis LSE_LINE_FILE_ID=38, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=78, LSE_RLINE=97 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(172[12] 188[10])
    defparam reg_04_i0_i31.GSR = "ENABLED";
    LUT4 wb_slave_data_31__I_0_i9_3_lut_4_lut (.A(write_ack_N_4033), .B(n41279), 
         .C(reg_00[8]), .D(wb_slave_data_31__N_3867[8]), .Z(\GPOwb_DAT_O[8] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(99[24] 100[31])
    defparam wb_slave_data_31__I_0_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 wb_slave_data_31__I_0_i2_3_lut_4_lut (.A(write_ack_N_4033), .B(n41279), 
         .C(GPOout_pins[1]), .D(wb_slave_data_31__N_3867[1]), .Z(\GPOwb_DAT_O[1] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(99[24] 100[31])
    defparam wb_slave_data_31__I_0_i2_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13368_3_lut_4_lut (.A(write_ack_N_4033), .B(n41279), .C(reg_00[16]), 
         .D(n18656), .Z(n13_adj_133)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(99[24] 100[31])
    defparam i13368_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13262_3_lut_4_lut (.A(write_ack_N_4033), .B(n41279), .C(reg_00[19]), 
         .D(n18553), .Z(n13_adj_134)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(99[24] 100[31])
    defparam i13262_3_lut_4_lut.init = 16'hfd20;
    LUT4 wb_slave_data_31__I_0_i1_4_lut (.A(n34304), .B(LED_G_c_0), .C(n41185), 
         .D(n34112), .Z(\GPOwb_DAT_O[0] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(114[23] 117[16])
    defparam wb_slave_data_31__I_0_i1_4_lut.init = 16'hcfca;
    LUT4 i13227_3_lut_4_lut (.A(write_ack_N_4033), .B(n41279), .C(reg_00[20]), 
         .D(n18519), .Z(n11)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(99[24] 100[31])
    defparam i13227_3_lut_4_lut.init = 16'hfd20;
    LUT4 i12980_3_lut_4_lut (.A(write_ack_N_4033), .B(n41279), .C(reg_00[27]), 
         .D(n18279), .Z(n13_adj_135)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(99[24] 100[31])
    defparam i12980_3_lut_4_lut.init = 16'hfd20;
    LUT4 wb_slave_data_31__I_0_i6_3_lut_4_lut (.A(write_ack_N_4033), .B(n41279), 
         .C(GPOout_pins[5]), .D(wb_slave_data_31__N_3867[5]), .Z(\GPOwb_DAT_O[5] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(99[24] 100[31])
    defparam wb_slave_data_31__I_0_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 i13508_3_lut_4_lut (.A(write_ack_N_4033), .B(n41279), .C(reg_00[12]), 
         .D(n18792), .Z(n13_adj_136)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(99[24] 100[31])
    defparam i13508_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5013_2_lut_3_lut_4_lut (.A(write_ack_N_4033), .B(n41279), .C(n41239), 
         .D(n41243), .Z(REF_CLK_c_enable_1511)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(99[24] 100[31])
    defparam i5013_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i4228_2_lut_3_lut_4_lut (.A(write_ack_N_4033), .B(n41279), .C(n41324), 
         .D(n41243), .Z(REF_CLK_c_enable_1487)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(99[24] 100[31])
    defparam i4228_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i4981_2_lut_3_lut_4_lut (.A(write_ack_N_4033), .B(n41279), .C(n41238), 
         .D(n41243), .Z(REF_CLK_c_enable_1495)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(99[24] 100[31])
    defparam i4981_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i12874_3_lut_4_lut (.A(write_ack_N_4033), .B(n41279), .C(reg_00[30]), 
         .D(n18176), .Z(n13_adj_137)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(99[24] 100[31])
    defparam i12874_3_lut_4_lut.init = 16'hfd20;
    LUT4 i30419_2_lut_rep_837 (.A(\SHAREDBUS_ADR_I[20] ), .B(\SHAREDBUS_ADR_I[29] ), 
         .Z(n41242)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i30419_2_lut_rep_837.init = 16'heeee;
    LUT4 i13362_3_lut_4_lut_4_lut (.A(write_ack_N_4033), .B(n41250), .C(reg_04_c[16]), 
         .D(n41251), .Z(n18656)) /* synthesis lut_function=((B (C+(D))+!B !((D)+!C))+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(103[24] 104[31])
    defparam i13362_3_lut_4_lut_4_lut.init = 16'hddf5;
    LUT4 i13256_3_lut_4_lut_4_lut (.A(write_ack_N_4033), .B(n41250), .C(reg_04_c[19]), 
         .D(n41251), .Z(n18553)) /* synthesis lut_function=((B (C+(D))+!B !((D)+!C))+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(103[24] 104[31])
    defparam i13256_3_lut_4_lut_4_lut.init = 16'hddf5;
    LUT4 i12974_3_lut_4_lut_4_lut (.A(write_ack_N_4033), .B(n41250), .C(reg_04_c[27]), 
         .D(n41251), .Z(n18279)) /* synthesis lut_function=((B (C+(D))+!B !((D)+!C))+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(103[24] 104[31])
    defparam i12974_3_lut_4_lut_4_lut.init = 16'hddf5;
    LUT4 i13115_3_lut_4_lut_4_lut (.A(write_ack_N_4033), .B(n41250), .C(reg_04_c[23]), 
         .D(n41251), .Z(n18416)) /* synthesis lut_function=((B (C+(D))+!B !((D)+!C))+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(103[24] 104[31])
    defparam i13115_3_lut_4_lut_4_lut.init = 16'hddf5;
    LUT4 i13010_3_lut_4_lut_4_lut (.A(write_ack_N_4033), .B(n41250), .C(reg_04_c[26]), 
         .D(n41251), .Z(n18314)) /* synthesis lut_function=((B (C+(D))+!B !((D)+!C))+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(103[24] 104[31])
    defparam i13010_3_lut_4_lut_4_lut.init = 16'hddf5;
    LUT4 wb_slave_data_31__I_166_i2_3_lut_4_lut_4_lut (.A(write_ack_N_4033), 
         .B(n41250), .C(reg_04_c[1]), .D(n41251), .Z(wb_slave_data_31__N_3867[1])) /* synthesis lut_function=((B (C+(D))+!B !((D)+!C))+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(103[24] 104[31])
    defparam wb_slave_data_31__I_166_i2_3_lut_4_lut_4_lut.init = 16'hddf5;
    LUT4 i1_4_lut_adj_260 (.A(n32388), .B(n41210), .C(n35914), .D(n35577), 
         .Z(write_ack_N_4033)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_260.init = 16'h0008;
    LUT4 i1_4_lut_adj_261 (.A(n15), .B(n35820), .C(n32366), .D(n41310), 
         .Z(n32388)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_261.init = 16'h0010;
    LUT4 i30752_4_lut (.A(n19), .B(n41225), .C(n35647), .D(n41258), 
         .Z(n35914)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30752_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_262 (.A(n35128), .B(n41210), .C(n15), .D(n35894), 
         .Z(write_ack_N_4031)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_262.init = 16'h0008;
    LUT4 i1_4_lut_adj_263 (.A(n35724), .B(n41225), .C(n19), .D(n35112), 
         .Z(n35128)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_263.init = 16'h0100;
    LUT4 i30732_4_lut (.A(n35647), .B(n41253), .C(n35583), .D(n41273), 
         .Z(n35894)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30732_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_264 (.A(n41243), .B(n41310), .C(n41246), .D(n41301), 
         .Z(n35112)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_4_lut_adj_264.init = 16'h2000;
    LUT4 i30439_2_lut (.A(\SHAREDBUS_ADR_I[26] ), .B(\SHAREDBUS_ADR_I[16] ), 
         .Z(n35583)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i30439_2_lut.init = 16'heeee;
    LUT4 i13572_3_lut_4_lut_4_lut (.A(write_ack_N_4033), .B(n41250), .C(reg_04_c[10]), 
         .D(n41251), .Z(n18860)) /* synthesis lut_function=((B (C+(D))+!B !((D)+!C))+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(103[24] 104[31])
    defparam i13572_3_lut_4_lut_4_lut.init = 16'hddf5;
    LUT4 i13221_3_lut_4_lut_4_lut (.A(write_ack_N_4033), .B(n41250), .C(reg_04_c[20]), 
         .D(n41251), .Z(n18519)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C+(D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(103[24] 104[31])
    defparam i13221_3_lut_4_lut_4_lut.init = 16'h22a0;
    LUT4 i13502_3_lut_4_lut_4_lut (.A(write_ack_N_4033), .B(n41250), .C(reg_04_c[12]), 
         .D(n41251), .Z(n18792)) /* synthesis lut_function=((B (C+(D))+!B !((D)+!C))+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(103[24] 104[31])
    defparam i13502_3_lut_4_lut_4_lut.init = 16'hddf5;
    LUT4 i12868_3_lut_4_lut_4_lut (.A(write_ack_N_4033), .B(n41250), .C(reg_04_c[30]), 
         .D(n41251), .Z(n18176)) /* synthesis lut_function=((B (C+(D))+!B !((D)+!C))+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(103[24] 104[31])
    defparam i12868_3_lut_4_lut_4_lut.init = 16'hddf5;
    LUT4 i12829_3_lut_4_lut_4_lut (.A(write_ack_N_4033), .B(n41250), .C(reg_04_c[31]), 
         .D(n41251), .Z(n18138)) /* synthesis lut_function=((B (C+(D))+!B !((D)+!C))+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(103[24] 104[31])
    defparam i12829_3_lut_4_lut_4_lut.init = 16'hddf5;
    LUT4 wb_slave_data_31__I_166_i9_3_lut_4_lut_4_lut (.A(write_ack_N_4033), 
         .B(n41250), .C(reg_04_c[8]), .D(n41251), .Z(wb_slave_data_31__N_3867[8])) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C+(D)))+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(103[24] 104[31])
    defparam wb_slave_data_31__I_166_i9_3_lut_4_lut_4_lut.init = 16'h22a0;
    LUT4 wb_slave_data_31__I_166_i6_3_lut_4_lut_4_lut (.A(write_ack_N_4033), 
         .B(n41250), .C(reg_04_c[5]), .D(n41251), .Z(wb_slave_data_31__N_3867[5])) /* synthesis lut_function=((B (C+(D))+!B !((D)+!C))+!A) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/Reg_Comp/rtl/verilog/wb_reg_dev.v(103[24] 104[31])
    defparam wb_slave_data_31__I_166_i6_3_lut_4_lut_4_lut.init = 16'hddf5;
    LUT4 i1_4_lut_adj_265 (.A(n35633), .B(n41210), .C(n32110), .D(n35898), 
         .Z(read_ack)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_adj_265.init = 16'h0040;
    LUT4 i1_4_lut_adj_266 (.A(n41269), .B(n41273), .C(n19), .D(n32096), 
         .Z(n32110)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_266.init = 16'h0100;
    LUT4 i30736_4_lut (.A(n41258), .B(n41260), .C(n34242), .D(n35739), 
         .Z(n35898)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30736_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_267 (.A(\SHAREDBUS_ADR_I[16] ), .B(n41304), .C(n41246), 
         .D(n41301), .Z(n32096)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_267.init = 16'h1000;
    LUT4 i1_4_lut_adj_268 (.A(n33318), .B(n35906), .C(n41225), .D(n19), 
         .Z(n33328)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_268.init = 16'h0002;
    LUT4 i1_4_lut_adj_269 (.A(n35577), .B(n41246), .C(n41310), .D(n33294), 
         .Z(n33318)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_269.init = 16'h0400;
    LUT4 i30744_4_lut (.A(n15), .B(n32312), .C(n35800), .D(n35583), 
         .Z(n35906)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30744_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_270 (.A(n33394), .B(n35906), .C(n41225), .D(n19), 
         .Z(n33404)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_270.init = 16'h0002;
    LUT4 i1_4_lut_adj_271 (.A(n35577), .B(n41246), .C(n41310), .D(n33370), 
         .Z(n33394)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_271.init = 16'h0400;
    LUT4 i1_4_lut_adj_272 (.A(n33280), .B(n35906), .C(n41225), .D(n19), 
         .Z(n33290)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_272.init = 16'h0002;
    LUT4 i30410_2_lut_rep_855 (.A(\SHAREDBUS_ADR_I[24] ), .B(\SHAREDBUS_ADR_I[25] ), 
         .Z(n41260)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i30410_2_lut_rep_855.init = 16'heeee;
    LUT4 i30425_2_lut_rep_868 (.A(\SHAREDBUS_ADR_I[18] ), .B(\SHAREDBUS_ADR_I[27] ), 
         .Z(n41273)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i30425_2_lut_rep_868.init = 16'heeee;
    LUT4 i30638_2_lut_3_lut_4_lut (.A(\SHAREDBUS_ADR_I[18] ), .B(\SHAREDBUS_ADR_I[27] ), 
         .C(\SHAREDBUS_ADR_I[29] ), .D(\SHAREDBUS_ADR_I[20] ), .Z(n35800)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30638_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i30658_2_lut_3_lut_4_lut (.A(\SHAREDBUS_ADR_I[18] ), .B(\SHAREDBUS_ADR_I[27] ), 
         .C(\SHAREDBUS_ADR_I[16] ), .D(\SHAREDBUS_ADR_I[22] ), .Z(n35820)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30658_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_273 (.A(n35577), .B(n41246), .C(n41310), .D(n33256), 
         .Z(n33280)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_273.init = 16'h0400;
    LUT4 i1_4_lut_adj_274 (.A(n33242), .B(n35906), .C(n41225), .D(n19), 
         .Z(n33252)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_274.init = 16'h0002;
    LUT4 i1_4_lut_adj_275 (.A(n35577), .B(n41246), .C(n41310), .D(n33218), 
         .Z(n33242)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_275.init = 16'h0400;
    LUT4 i1_4_lut_adj_276 (.A(n33204), .B(n35906), .C(n41225), .D(n19), 
         .Z(n33214)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_276.init = 16'h0002;
    LUT4 i1_4_lut_adj_277 (.A(n35577), .B(n41246), .C(n41310), .D(n33180), 
         .Z(n33204)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_277.init = 16'h0400;
    LUT4 i1_4_lut_adj_278 (.A(n33356), .B(n35906), .C(n41225), .D(n19), 
         .Z(n33366)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_278.init = 16'h0002;
    
endmodule
//
// Verilog Description of module \gpio(DATA_WIDTH=32'b01,INPUT_WIDTH=32'b01,OUTPUT_WIDTH=32'b01,EDGE=1,POSE_EDGE_IRQ=1,INPUT_PORTS_ONLY=0,BOTH_INPUT_AND_OUTPUT=1) 
//

module \gpio(DATA_WIDTH=32'b01,INPUT_WIDTH=32'b01,OUTPUT_WIDTH=32'b01,EDGE=1,POSE_EDGE_IRQ=1,INPUT_PORTS_ONLY=0,BOTH_INPUT_AND_OUTPUT=1)  (GPIOGPIO_ACK_O, 
            REF_CLK_c, REF_CLK_c_enable_1606, PIO_DATAI_0__N_3822, LED_B_c_0, 
            REF_CLK_c_enable_424, n36339, PIO_DATAI, n36340, n35006, 
            PIO_OUT_7__N_3493, n41275, n41310, \SHAREDBUS_ADR_I[7] , 
            n954, LEDGPIO_ACK_O) /* synthesis syn_module_defined=1 */ ;
    output GPIOGPIO_ACK_O;
    input REF_CLK_c;
    input REF_CLK_c_enable_1606;
    input PIO_DATAI_0__N_3822;
    output LED_B_c_0;
    input REF_CLK_c_enable_424;
    input n36339;
    output [0:0]PIO_DATAI;
    input n36340;
    output n35006;
    output PIO_OUT_7__N_3493;
    input n41275;
    input n41310;
    input \SHAREDBUS_ADR_I[7] ;
    input [0:0]n954;
    input LEDGPIO_ACK_O;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    
    wire n34998;
    
    FD1S3DX GPIO_ACK_O_108 (.D(PIO_DATAI_0__N_3822), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(GPIOGPIO_ACK_O)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=707, LSE_RLINE=724 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/gpio/rtl/verilog/gpio.v(188[11] 191[33])
    defparam GPIO_ACK_O_108.GSR = "ENABLED";
    FD1P3DX PIO_DATAO_0__109 (.D(n36339), .SP(REF_CLK_c_enable_424), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(LED_B_c_0)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=707, LSE_RLINE=724 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/gpio/rtl/verilog/gpio.v(396[11] 397[65])
    defparam PIO_DATAO_0__109.GSR = "ENABLED";
    FD1P3DX PIO_DATAI_0__110 (.D(n36340), .SP(REF_CLK_c_enable_424), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(PIO_DATAI[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=707, LSE_RLINE=724 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/gpio/rtl/verilog/gpio.v(438[11] 439[59])
    defparam PIO_DATAI_0__110.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(n35006), .B(REF_CLK_c_enable_424), .Z(PIO_OUT_7__N_3493)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_4_lut (.A(n41275), .B(n41310), .C(\SHAREDBUS_ADR_I[7] ), .D(n34998), 
         .Z(n35006)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_adj_259 (.A(n954[0]), .B(LEDGPIO_ACK_O), .Z(n34998)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_259.init = 16'h2222;
    
endmodule
//
// Verilog Description of module \FIFO_Comp(reg_16_int_val=32'b010010001101001010101111001101) 
//

module \FIFO_Comp(reg_16_int_val=32'b010010001101001010101111001101)  (n32828, 
            n41246, n34372, n5223, n15, n41303, \SHAREDBUS_ADR_I[25] , 
            \SHAREDBUS_ADR_I[24] , \SHAREDBUS_ADR_I[29] , \SHAREDBUS_ADR_I[16] , 
            n41345, \SHAREDBUS_ADR_I[7] , n41186, n16, n17, n19, 
            n5, read_ack, REF_CLK_c, REF_CLK_c_enable_1606, n31476, 
            n19_adj_66, n5_adj_67, n16_adj_68, n17_adj_69, n16_adj_70, 
            n22, n16_adj_71, n22_adj_72, n8, n2, n16_adj_73, n22_adj_74, 
            n16_adj_75, n22_adj_76, n8_adj_77, n2_adj_78, n41344, 
            n19_adj_79, n26, n359, n392, n16_adj_80, n17_adj_81, 
            n16_adj_82, n17_adj_83, n17_adj_84, n5_adj_85, n13, n14, 
            REF_CLK_c_enable_1550, n41328, inst1_FIFOfifo_rst, REF_CLK_c_enable_1581, 
            write_ack, write_ack_N_4649, inst3_Empty, fiford_reg, fiford, 
            n40677, \SHAREDBUS_ADR_I[23] , \SHAREDBUS_ADR_I[18] , n32798, 
            inst3_Q, n41347, n31779, n41329, n41330, n41331, n41332, 
            n41333, n41334, n41335, REF_CLK_c_enable_1558, \SHAREDBUS_DAT_I[8] , 
            \SHAREDBUS_DAT_I[9] , \SHAREDBUS_DAT_I[10] , \SHAREDBUS_DAT_I[11] , 
            \SHAREDBUS_DAT_I[12] , \SHAREDBUS_DAT_I[13] , \SHAREDBUS_DAT_I[14] , 
            \SHAREDBUS_DAT_I[15] , REF_CLK_c_enable_1566, n41336, n41337, 
            n41338, n41339, n41340, n41341, n41342, n41343, REF_CLK_c_enable_1574, 
            \SHAREDBUS_DAT_I[24] , \SHAREDBUS_DAT_I[25] , \SHAREDBUS_DAT_I[26] , 
            \SHAREDBUS_DAT_I[27] , \SHAREDBUS_DAT_I[28] , \SHAREDBUS_DAT_I[29] , 
            \SHAREDBUS_DAT_I[30] , \SHAREDBUS_DAT_I[31] , \reg_12[2] , 
            \reg_12[3] , \reg_12[4] , \reg_12[6] , \reg_12[7] , REF_CLK_c_enable_1589, 
            \reg_12[9] , \reg_12[11] , \reg_12[12] , \reg_12[13] , \reg_12[14] , 
            \reg_12[15] , REF_CLK_c_enable_1597, \reg_12[17] , \reg_12[18] , 
            \reg_12[21] , \reg_12[22] , \reg_12[24] , REF_CLK_c_enable_1605, 
            \reg_12[25] , \reg_12[28] , \reg_12[29] , inst3_Full, n41193, 
            n2_adj_86, n37903, n2_adj_87, n37905, n2_adj_88, n4893, 
            n2_adj_89, n2_adj_90, n2_adj_91, n2_adj_92, n37904, n2_adj_93, 
            n2_adj_94, n4883, n2_adj_95, n2_adj_96, n4880, n2_adj_97, 
            n2_adj_98, n37906, n2_adj_99, n4875, n2_adj_100, n4873, 
            n2_adj_101, n41275, REF_CLK_c_enable_424, n41310, n30762, 
            n30241, n41180, n41181, \FIFOwb_DAT_O[12] , n2_adj_102, 
            n2_adj_103, n4868, n954, n953, n41301, n32366, n41262, 
            n41278, n35136, n33088, n41304, n34742, n41226, n41255, 
            n41323, n5_adj_104, spiSPI_ACK_O, n35042, n352, n385, 
            n19_adj_105, n26_adj_106, n19_adj_107, n25, n19_adj_108, 
            n25_adj_109, n355, n388, n19_adj_110, n5_adj_111, n19_adj_112, 
            n25_adj_113, n17_adj_114, n22_adj_115, n8_adj_116, n2_adj_117, 
            n19_adj_118, n25_adj_119, n19_adj_120, n25_adj_121, n360, 
            n393, n31183, n23, n31, n19_adj_122, n5_adj_123, n8_adj_124, 
            n2_adj_125, n19_adj_126, n25_adj_127, n19_adj_128, n5_adj_129, 
            n33846, \FIFOwb_DAT_O[0] , n41210, n33864, n19_adj_130, 
            n41258, n30949, \SHAREDBUS_ADR_I[30] , n41272, n41265, 
            n30951, n30948, n30944, \SHAREDBUS_ADR_I[20] , \SHAREDBUS_ADR_I[26] , 
            \SHAREDBUS_ADR_I[27] , \SHAREDBUS_ADR_I[22] , n35844, n35866, 
            n41274, \SHAREDBUS_ADR_I[5] , n41346, n41225, n35633, 
            n35736, n41277, n41289, n32814, n35796, \FIFOwb_DAT_O[18] , 
            \FIFOwb_DAT_O[25] , n37954, \FIFOwb_DAT_O[31] , n37956, 
            \FIFOwb_DAT_O[30] , n37955, \FIFOwb_DAT_O[27] , \FIFOwb_DAT_O[26] , 
            \FIFOwb_DAT_O[23] , \FIFOwb_DAT_O[20] , \FIFOwb_DAT_O[19] , 
            \FIFOwb_DAT_O[16] , \FIFOwb_DAT_O[10] , \FIFOwb_DAT_O[8] , 
            \FIFOwb_DAT_O[5] , \FIFOwb_DAT_O[1] , \FIFOwb_DAT_O[21] , 
            \FIFOwb_DAT_O[28] , \FIFOwb_DAT_O[15] , \FIFOwb_DAT_O[13] , 
            \FIFOwb_DAT_O[11] , \FIFOwb_DAT_O[9] ) /* synthesis syn_module_defined=1 */ ;
    input n32828;
    output n41246;
    output n34372;
    output n5223;
    input n15;
    input n41303;
    input \SHAREDBUS_ADR_I[25] ;
    input \SHAREDBUS_ADR_I[24] ;
    input \SHAREDBUS_ADR_I[29] ;
    input \SHAREDBUS_ADR_I[16] ;
    input n41345;
    input \SHAREDBUS_ADR_I[7] ;
    output n41186;
    input n16;
    output n17;
    input n19;
    output n5;
    output read_ack;
    input REF_CLK_c;
    input REF_CLK_c_enable_1606;
    input n31476;
    input n19_adj_66;
    output n5_adj_67;
    input n16_adj_68;
    output n17_adj_69;
    input n16_adj_70;
    output n22;
    input n16_adj_71;
    output n22_adj_72;
    input n8;
    output n2;
    input n16_adj_73;
    output n22_adj_74;
    input n16_adj_75;
    output n22_adj_76;
    input n8_adj_77;
    output n2_adj_78;
    input n41344;
    input n19_adj_79;
    output n26;
    input n359;
    output n392;
    input n16_adj_80;
    output n17_adj_81;
    input n16_adj_82;
    output n17_adj_83;
    input n17_adj_84;
    output n5_adj_85;
    input n13;
    output n14;
    input REF_CLK_c_enable_1550;
    input n41328;
    output inst1_FIFOfifo_rst;
    input REF_CLK_c_enable_1581;
    output write_ack;
    input write_ack_N_4649;
    input inst3_Empty;
    output fiford_reg;
    input fiford;
    input n40677;
    input \SHAREDBUS_ADR_I[23] ;
    input \SHAREDBUS_ADR_I[18] ;
    output n32798;
    input [31:0]inst3_Q;
    input n41347;
    output n31779;
    input n41329;
    input n41330;
    input n41331;
    input n41332;
    input n41333;
    input n41334;
    input n41335;
    input REF_CLK_c_enable_1558;
    input \SHAREDBUS_DAT_I[8] ;
    input \SHAREDBUS_DAT_I[9] ;
    input \SHAREDBUS_DAT_I[10] ;
    input \SHAREDBUS_DAT_I[11] ;
    input \SHAREDBUS_DAT_I[12] ;
    input \SHAREDBUS_DAT_I[13] ;
    input \SHAREDBUS_DAT_I[14] ;
    input \SHAREDBUS_DAT_I[15] ;
    input REF_CLK_c_enable_1566;
    input n41336;
    input n41337;
    input n41338;
    input n41339;
    input n41340;
    input n41341;
    input n41342;
    input n41343;
    input REF_CLK_c_enable_1574;
    input \SHAREDBUS_DAT_I[24] ;
    input \SHAREDBUS_DAT_I[25] ;
    input \SHAREDBUS_DAT_I[26] ;
    input \SHAREDBUS_DAT_I[27] ;
    input \SHAREDBUS_DAT_I[28] ;
    input \SHAREDBUS_DAT_I[29] ;
    input \SHAREDBUS_DAT_I[30] ;
    input \SHAREDBUS_DAT_I[31] ;
    output \reg_12[2] ;
    output \reg_12[3] ;
    output \reg_12[4] ;
    output \reg_12[6] ;
    output \reg_12[7] ;
    input REF_CLK_c_enable_1589;
    output \reg_12[9] ;
    output \reg_12[11] ;
    output \reg_12[12] ;
    output \reg_12[13] ;
    output \reg_12[14] ;
    output \reg_12[15] ;
    input REF_CLK_c_enable_1597;
    output \reg_12[17] ;
    output \reg_12[18] ;
    output \reg_12[21] ;
    output \reg_12[22] ;
    output \reg_12[24] ;
    input REF_CLK_c_enable_1605;
    output \reg_12[25] ;
    output \reg_12[28] ;
    output \reg_12[29] ;
    input inst3_Full;
    input n41193;
    input n2_adj_86;
    input n37903;
    input n2_adj_87;
    input n37905;
    input n2_adj_88;
    output n4893;
    input n2_adj_89;
    input n2_adj_90;
    input n2_adj_91;
    input n2_adj_92;
    input n37904;
    input n2_adj_93;
    input n2_adj_94;
    output n4883;
    input n2_adj_95;
    input n2_adj_96;
    output n4880;
    input n2_adj_97;
    input n2_adj_98;
    input n37906;
    input n2_adj_99;
    output n4875;
    input n2_adj_100;
    output n4873;
    input n2_adj_101;
    input n41275;
    input REF_CLK_c_enable_424;
    input n41310;
    input n30762;
    output n30241;
    output n41180;
    output n41181;
    output \FIFOwb_DAT_O[12] ;
    input n2_adj_102;
    input n2_adj_103;
    output n4868;
    input [0:0]n954;
    input [0:0]n953;
    input n41301;
    output n32366;
    input n41262;
    input n41278;
    output n35136;
    output n33088;
    input n41304;
    output n34742;
    output n41226;
    input n41255;
    input n41323;
    output n5_adj_104;
    input spiSPI_ACK_O;
    output n35042;
    input n352;
    output n385;
    input n19_adj_105;
    output n26_adj_106;
    input n19_adj_107;
    output n25;
    input n19_adj_108;
    output n25_adj_109;
    input n355;
    output n388;
    input n19_adj_110;
    output n5_adj_111;
    input n19_adj_112;
    output n25_adj_113;
    input n17_adj_114;
    output n22_adj_115;
    input n8_adj_116;
    output n2_adj_117;
    input n19_adj_118;
    output n25_adj_119;
    input n19_adj_120;
    output n25_adj_121;
    input n360;
    output n393;
    input n31183;
    input n23;
    output n31;
    input n19_adj_122;
    output n5_adj_123;
    input n8_adj_124;
    output n2_adj_125;
    input n19_adj_126;
    output n25_adj_127;
    input n19_adj_128;
    output n5_adj_129;
    output n33846;
    output \FIFOwb_DAT_O[0] ;
    input n41210;
    input n33864;
    input n19_adj_130;
    output n41258;
    output n30949;
    input \SHAREDBUS_ADR_I[30] ;
    output n41272;
    input n41265;
    output n30951;
    output n30948;
    output n30944;
    input \SHAREDBUS_ADR_I[20] ;
    input \SHAREDBUS_ADR_I[26] ;
    input \SHAREDBUS_ADR_I[27] ;
    input \SHAREDBUS_ADR_I[22] ;
    output n35844;
    output n35866;
    output n41274;
    input \SHAREDBUS_ADR_I[5] ;
    input n41346;
    output n41225;
    output n35633;
    output n35736;
    output n41277;
    input n41289;
    output n32814;
    output n35796;
    output \FIFOwb_DAT_O[18] ;
    output \FIFOwb_DAT_O[25] ;
    input n37954;
    output \FIFOwb_DAT_O[31] ;
    input n37956;
    output \FIFOwb_DAT_O[30] ;
    input n37955;
    output \FIFOwb_DAT_O[27] ;
    output \FIFOwb_DAT_O[26] ;
    output \FIFOwb_DAT_O[23] ;
    output \FIFOwb_DAT_O[20] ;
    output \FIFOwb_DAT_O[19] ;
    output \FIFOwb_DAT_O[16] ;
    output \FIFOwb_DAT_O[10] ;
    output \FIFOwb_DAT_O[8] ;
    output \FIFOwb_DAT_O[5] ;
    output \FIFOwb_DAT_O[1] ;
    output \FIFOwb_DAT_O[21] ;
    output \FIFOwb_DAT_O[28] ;
    output \FIFOwb_DAT_O[15] ;
    output \FIFOwb_DAT_O[13] ;
    output \FIFOwb_DAT_O[11] ;
    output \FIFOwb_DAT_O[9] ;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    
    wb_fifo_dev instantiate_wb_fifo_dev (.n32828(n32828), .n41246(n41246), 
            .n34372(n34372), .n5223(n5223), .n15(n15), .n41303(n41303), 
            .\SHAREDBUS_ADR_I[25] (\SHAREDBUS_ADR_I[25] ), .\SHAREDBUS_ADR_I[24] (\SHAREDBUS_ADR_I[24] ), 
            .\SHAREDBUS_ADR_I[29] (\SHAREDBUS_ADR_I[29] ), .\SHAREDBUS_ADR_I[16] (\SHAREDBUS_ADR_I[16] ), 
            .n41345(n41345), .\SHAREDBUS_ADR_I[7] (\SHAREDBUS_ADR_I[7] ), 
            .n41186(n41186), .n16(n16), .n17(n17), .n19(n19), .n5(n5), 
            .read_ack(read_ack), .REF_CLK_c(REF_CLK_c), .REF_CLK_c_enable_1606(REF_CLK_c_enable_1606), 
            .n31476(n31476), .n19_adj_1(n19_adj_66), .n5_adj_2(n5_adj_67), 
            .n16_adj_3(n16_adj_68), .n17_adj_4(n17_adj_69), .n16_adj_5(n16_adj_70), 
            .n22(n22), .n16_adj_6(n16_adj_71), .n22_adj_7(n22_adj_72), 
            .n8(n8), .n2(n2), .n16_adj_8(n16_adj_73), .n22_adj_9(n22_adj_74), 
            .n16_adj_10(n16_adj_75), .n22_adj_11(n22_adj_76), .n8_adj_12(n8_adj_77), 
            .n2_adj_13(n2_adj_78), .n41344(n41344), .n19_adj_14(n19_adj_79), 
            .n26(n26), .n359(n359), .n392(n392), .n16_adj_15(n16_adj_80), 
            .n17_adj_16(n17_adj_81), .n16_adj_17(n16_adj_82), .n17_adj_18(n17_adj_83), 
            .n17_adj_19(n17_adj_84), .n5_adj_20(n5_adj_85), .n13(n13), 
            .n14(n14), .REF_CLK_c_enable_1550(REF_CLK_c_enable_1550), .n41328(n41328), 
            .inst1_FIFOfifo_rst(inst1_FIFOfifo_rst), .REF_CLK_c_enable_1581(REF_CLK_c_enable_1581), 
            .write_ack(write_ack), .write_ack_N_4649(write_ack_N_4649), 
            .inst3_Empty(inst3_Empty), .fiford_reg(fiford_reg), .fiford(fiford), 
            .n40677(n40677), .\SHAREDBUS_ADR_I[23] (\SHAREDBUS_ADR_I[23] ), 
            .\SHAREDBUS_ADR_I[18] (\SHAREDBUS_ADR_I[18] ), .n32798(n32798), 
            .inst3_Q({inst3_Q}), .n41347(n41347), .n31779(n31779), .n41329(n41329), 
            .n41330(n41330), .n41331(n41331), .n41332(n41332), .n41333(n41333), 
            .n41334(n41334), .n41335(n41335), .REF_CLK_c_enable_1558(REF_CLK_c_enable_1558), 
            .\SHAREDBUS_DAT_I[8] (\SHAREDBUS_DAT_I[8] ), .\SHAREDBUS_DAT_I[9] (\SHAREDBUS_DAT_I[9] ), 
            .\SHAREDBUS_DAT_I[10] (\SHAREDBUS_DAT_I[10] ), .\SHAREDBUS_DAT_I[11] (\SHAREDBUS_DAT_I[11] ), 
            .\SHAREDBUS_DAT_I[12] (\SHAREDBUS_DAT_I[12] ), .\SHAREDBUS_DAT_I[13] (\SHAREDBUS_DAT_I[13] ), 
            .\SHAREDBUS_DAT_I[14] (\SHAREDBUS_DAT_I[14] ), .\SHAREDBUS_DAT_I[15] (\SHAREDBUS_DAT_I[15] ), 
            .REF_CLK_c_enable_1566(REF_CLK_c_enable_1566), .n41336(n41336), 
            .n41337(n41337), .n41338(n41338), .n41339(n41339), .n41340(n41340), 
            .n41341(n41341), .n41342(n41342), .n41343(n41343), .REF_CLK_c_enable_1574(REF_CLK_c_enable_1574), 
            .\SHAREDBUS_DAT_I[24] (\SHAREDBUS_DAT_I[24] ), .\SHAREDBUS_DAT_I[25] (\SHAREDBUS_DAT_I[25] ), 
            .\SHAREDBUS_DAT_I[26] (\SHAREDBUS_DAT_I[26] ), .\SHAREDBUS_DAT_I[27] (\SHAREDBUS_DAT_I[27] ), 
            .\SHAREDBUS_DAT_I[28] (\SHAREDBUS_DAT_I[28] ), .\SHAREDBUS_DAT_I[29] (\SHAREDBUS_DAT_I[29] ), 
            .\SHAREDBUS_DAT_I[30] (\SHAREDBUS_DAT_I[30] ), .\SHAREDBUS_DAT_I[31] (\SHAREDBUS_DAT_I[31] ), 
            .\reg_12[2] (\reg_12[2] ), .\reg_12[3] (\reg_12[3] ), .\reg_12[4] (\reg_12[4] ), 
            .\reg_12[6] (\reg_12[6] ), .\reg_12[7] (\reg_12[7] ), .REF_CLK_c_enable_1589(REF_CLK_c_enable_1589), 
            .\reg_12[9] (\reg_12[9] ), .\reg_12[11] (\reg_12[11] ), .\reg_12[12] (\reg_12[12] ), 
            .\reg_12[13] (\reg_12[13] ), .\reg_12[14] (\reg_12[14] ), .\reg_12[15] (\reg_12[15] ), 
            .REF_CLK_c_enable_1597(REF_CLK_c_enable_1597), .\reg_12[17] (\reg_12[17] ), 
            .\reg_12[18] (\reg_12[18] ), .\reg_12[21] (\reg_12[21] ), .\reg_12[22] (\reg_12[22] ), 
            .\reg_12[24] (\reg_12[24] ), .REF_CLK_c_enable_1605(REF_CLK_c_enable_1605), 
            .\reg_12[25] (\reg_12[25] ), .\reg_12[28] (\reg_12[28] ), .\reg_12[29] (\reg_12[29] ), 
            .inst3_Full(inst3_Full), .n41193(n41193), .n2_adj_21(n2_adj_86), 
            .n37903(n37903), .n2_adj_22(n2_adj_87), .n37905(n37905), .n2_adj_23(n2_adj_88), 
            .n4893(n4893), .n2_adj_24(n2_adj_89), .n2_adj_25(n2_adj_90), 
            .n2_adj_26(n2_adj_91), .n2_adj_27(n2_adj_92), .n37904(n37904), 
            .n2_adj_28(n2_adj_93), .n2_adj_29(n2_adj_94), .n4883(n4883), 
            .n2_adj_30(n2_adj_95), .n2_adj_31(n2_adj_96), .n4880(n4880), 
            .n2_adj_32(n2_adj_97), .n2_adj_33(n2_adj_98), .n37906(n37906), 
            .n2_adj_34(n2_adj_99), .n4875(n4875), .n2_adj_35(n2_adj_100), 
            .n4873(n4873), .n2_adj_36(n2_adj_101), .n41275(n41275), .REF_CLK_c_enable_424(REF_CLK_c_enable_424), 
            .n41310(n41310), .n30762(n30762), .n30241(n30241), .n41180(n41180), 
            .n41181(n41181), .\FIFOwb_DAT_O[12] (\FIFOwb_DAT_O[12] ), .n2_adj_37(n2_adj_102), 
            .n2_adj_38(n2_adj_103), .n4868(n4868), .n954({n954}), .n953({n953}), 
            .n41301(n41301), .n32366(n32366), .n41262(n41262), .n41278(n41278), 
            .n35136(n35136), .n33088(n33088), .n41304(n41304), .n34742(n34742), 
            .n41226(n41226), .n41255(n41255), .n41323(n41323), .n5_adj_39(n5_adj_104), 
            .spiSPI_ACK_O(spiSPI_ACK_O), .n35042(n35042), .n352(n352), 
            .n385(n385), .n19_adj_40(n19_adj_105), .n26_adj_41(n26_adj_106), 
            .n19_adj_42(n19_adj_107), .n25(n25), .n19_adj_43(n19_adj_108), 
            .n25_adj_44(n25_adj_109), .n355(n355), .n388(n388), .n19_adj_45(n19_adj_110), 
            .n5_adj_46(n5_adj_111), .n19_adj_47(n19_adj_112), .n25_adj_48(n25_adj_113), 
            .n17_adj_49(n17_adj_114), .n22_adj_50(n22_adj_115), .n8_adj_51(n8_adj_116), 
            .n2_adj_52(n2_adj_117), .n19_adj_53(n19_adj_118), .n25_adj_54(n25_adj_119), 
            .n19_adj_55(n19_adj_120), .n25_adj_56(n25_adj_121), .n360(n360), 
            .n393(n393), .n31183(n31183), .n23(n23), .n31(n31), .n19_adj_57(n19_adj_122), 
            .n5_adj_58(n5_adj_123), .n8_adj_59(n8_adj_124), .n2_adj_60(n2_adj_125), 
            .n19_adj_61(n19_adj_126), .n25_adj_62(n25_adj_127), .n19_adj_63(n19_adj_128), 
            .n5_adj_64(n5_adj_129), .n33846(n33846), .\FIFOwb_DAT_O[0] (\FIFOwb_DAT_O[0] ), 
            .n41210(n41210), .n33864(n33864), .n19_adj_65(n19_adj_130), 
            .n41258(n41258), .n30949(n30949), .\SHAREDBUS_ADR_I[30] (\SHAREDBUS_ADR_I[30] ), 
            .n41272(n41272), .n41265(n41265), .n30951(n30951), .n30948(n30948), 
            .n30944(n30944), .\SHAREDBUS_ADR_I[20] (\SHAREDBUS_ADR_I[20] ), 
            .\SHAREDBUS_ADR_I[26] (\SHAREDBUS_ADR_I[26] ), .\SHAREDBUS_ADR_I[27] (\SHAREDBUS_ADR_I[27] ), 
            .\SHAREDBUS_ADR_I[22] (\SHAREDBUS_ADR_I[22] ), .n35844(n35844), 
            .n35866(n35866), .n41274(n41274), .\SHAREDBUS_ADR_I[5] (\SHAREDBUS_ADR_I[5] ), 
            .n41346(n41346), .n41225(n41225), .n35633(n35633), .n35736(n35736), 
            .n41277(n41277), .n41289(n41289), .n32814(n32814), .n35796(n35796), 
            .\FIFOwb_DAT_O[18] (\FIFOwb_DAT_O[18] ), .\FIFOwb_DAT_O[25] (\FIFOwb_DAT_O[25] ), 
            .n37954(n37954), .\FIFOwb_DAT_O[31] (\FIFOwb_DAT_O[31] ), .n37956(n37956), 
            .\FIFOwb_DAT_O[30] (\FIFOwb_DAT_O[30] ), .n37955(n37955), .\FIFOwb_DAT_O[27] (\FIFOwb_DAT_O[27] ), 
            .\FIFOwb_DAT_O[26] (\FIFOwb_DAT_O[26] ), .\FIFOwb_DAT_O[23] (\FIFOwb_DAT_O[23] ), 
            .\FIFOwb_DAT_O[20] (\FIFOwb_DAT_O[20] ), .\FIFOwb_DAT_O[19] (\FIFOwb_DAT_O[19] ), 
            .\FIFOwb_DAT_O[16] (\FIFOwb_DAT_O[16] ), .\FIFOwb_DAT_O[10] (\FIFOwb_DAT_O[10] ), 
            .\FIFOwb_DAT_O[8] (\FIFOwb_DAT_O[8] ), .\FIFOwb_DAT_O[5] (\FIFOwb_DAT_O[5] ), 
            .\FIFOwb_DAT_O[1] (\FIFOwb_DAT_O[1] ), .\FIFOwb_DAT_O[21] (\FIFOwb_DAT_O[21] ), 
            .\FIFOwb_DAT_O[28] (\FIFOwb_DAT_O[28] ), .\FIFOwb_DAT_O[15] (\FIFOwb_DAT_O[15] ), 
            .\FIFOwb_DAT_O[13] (\FIFOwb_DAT_O[13] ), .\FIFOwb_DAT_O[11] (\FIFOwb_DAT_O[11] ), 
            .\FIFOwb_DAT_O[9] (\FIFOwb_DAT_O[9] )) /* synthesis syn_module_defined=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/FIFO_Comp.v(83[11] 109[34])
    
endmodule
//
// Verilog Description of module wb_fifo_dev
//

module wb_fifo_dev (n32828, n41246, n34372, n5223, n15, n41303, 
            \SHAREDBUS_ADR_I[25] , \SHAREDBUS_ADR_I[24] , \SHAREDBUS_ADR_I[29] , 
            \SHAREDBUS_ADR_I[16] , n41345, \SHAREDBUS_ADR_I[7] , n41186, 
            n16, n17, n19, n5, read_ack, REF_CLK_c, REF_CLK_c_enable_1606, 
            n31476, n19_adj_1, n5_adj_2, n16_adj_3, n17_adj_4, n16_adj_5, 
            n22, n16_adj_6, n22_adj_7, n8, n2, n16_adj_8, n22_adj_9, 
            n16_adj_10, n22_adj_11, n8_adj_12, n2_adj_13, n41344, 
            n19_adj_14, n26, n359, n392, n16_adj_15, n17_adj_16, 
            n16_adj_17, n17_adj_18, n17_adj_19, n5_adj_20, n13, n14, 
            REF_CLK_c_enable_1550, n41328, inst1_FIFOfifo_rst, REF_CLK_c_enable_1581, 
            write_ack, write_ack_N_4649, inst3_Empty, fiford_reg, fiford, 
            n40677, \SHAREDBUS_ADR_I[23] , \SHAREDBUS_ADR_I[18] , n32798, 
            inst3_Q, n41347, n31779, n41329, n41330, n41331, n41332, 
            n41333, n41334, n41335, REF_CLK_c_enable_1558, \SHAREDBUS_DAT_I[8] , 
            \SHAREDBUS_DAT_I[9] , \SHAREDBUS_DAT_I[10] , \SHAREDBUS_DAT_I[11] , 
            \SHAREDBUS_DAT_I[12] , \SHAREDBUS_DAT_I[13] , \SHAREDBUS_DAT_I[14] , 
            \SHAREDBUS_DAT_I[15] , REF_CLK_c_enable_1566, n41336, n41337, 
            n41338, n41339, n41340, n41341, n41342, n41343, REF_CLK_c_enable_1574, 
            \SHAREDBUS_DAT_I[24] , \SHAREDBUS_DAT_I[25] , \SHAREDBUS_DAT_I[26] , 
            \SHAREDBUS_DAT_I[27] , \SHAREDBUS_DAT_I[28] , \SHAREDBUS_DAT_I[29] , 
            \SHAREDBUS_DAT_I[30] , \SHAREDBUS_DAT_I[31] , \reg_12[2] , 
            \reg_12[3] , \reg_12[4] , \reg_12[6] , \reg_12[7] , REF_CLK_c_enable_1589, 
            \reg_12[9] , \reg_12[11] , \reg_12[12] , \reg_12[13] , \reg_12[14] , 
            \reg_12[15] , REF_CLK_c_enable_1597, \reg_12[17] , \reg_12[18] , 
            \reg_12[21] , \reg_12[22] , \reg_12[24] , REF_CLK_c_enable_1605, 
            \reg_12[25] , \reg_12[28] , \reg_12[29] , inst3_Full, n41193, 
            n2_adj_21, n37903, n2_adj_22, n37905, n2_adj_23, n4893, 
            n2_adj_24, n2_adj_25, n2_adj_26, n2_adj_27, n37904, n2_adj_28, 
            n2_adj_29, n4883, n2_adj_30, n2_adj_31, n4880, n2_adj_32, 
            n2_adj_33, n37906, n2_adj_34, n4875, n2_adj_35, n4873, 
            n2_adj_36, n41275, REF_CLK_c_enable_424, n41310, n30762, 
            n30241, n41180, n41181, \FIFOwb_DAT_O[12] , n2_adj_37, 
            n2_adj_38, n4868, n954, n953, n41301, n32366, n41262, 
            n41278, n35136, n33088, n41304, n34742, n41226, n41255, 
            n41323, n5_adj_39, spiSPI_ACK_O, n35042, n352, n385, 
            n19_adj_40, n26_adj_41, n19_adj_42, n25, n19_adj_43, n25_adj_44, 
            n355, n388, n19_adj_45, n5_adj_46, n19_adj_47, n25_adj_48, 
            n17_adj_49, n22_adj_50, n8_adj_51, n2_adj_52, n19_adj_53, 
            n25_adj_54, n19_adj_55, n25_adj_56, n360, n393, n31183, 
            n23, n31, n19_adj_57, n5_adj_58, n8_adj_59, n2_adj_60, 
            n19_adj_61, n25_adj_62, n19_adj_63, n5_adj_64, n33846, 
            \FIFOwb_DAT_O[0] , n41210, n33864, n19_adj_65, n41258, 
            n30949, \SHAREDBUS_ADR_I[30] , n41272, n41265, n30951, 
            n30948, n30944, \SHAREDBUS_ADR_I[20] , \SHAREDBUS_ADR_I[26] , 
            \SHAREDBUS_ADR_I[27] , \SHAREDBUS_ADR_I[22] , n35844, n35866, 
            n41274, \SHAREDBUS_ADR_I[5] , n41346, n41225, n35633, 
            n35736, n41277, n41289, n32814, n35796, \FIFOwb_DAT_O[18] , 
            \FIFOwb_DAT_O[25] , n37954, \FIFOwb_DAT_O[31] , n37956, 
            \FIFOwb_DAT_O[30] , n37955, \FIFOwb_DAT_O[27] , \FIFOwb_DAT_O[26] , 
            \FIFOwb_DAT_O[23] , \FIFOwb_DAT_O[20] , \FIFOwb_DAT_O[19] , 
            \FIFOwb_DAT_O[16] , \FIFOwb_DAT_O[10] , \FIFOwb_DAT_O[8] , 
            \FIFOwb_DAT_O[5] , \FIFOwb_DAT_O[1] , \FIFOwb_DAT_O[21] , 
            \FIFOwb_DAT_O[28] , \FIFOwb_DAT_O[15] , \FIFOwb_DAT_O[13] , 
            \FIFOwb_DAT_O[11] , \FIFOwb_DAT_O[9] ) /* synthesis syn_module_defined=1 */ ;
    input n32828;
    output n41246;
    output n34372;
    output n5223;
    input n15;
    input n41303;
    input \SHAREDBUS_ADR_I[25] ;
    input \SHAREDBUS_ADR_I[24] ;
    input \SHAREDBUS_ADR_I[29] ;
    input \SHAREDBUS_ADR_I[16] ;
    input n41345;
    input \SHAREDBUS_ADR_I[7] ;
    output n41186;
    input n16;
    output n17;
    input n19;
    output n5;
    output read_ack;
    input REF_CLK_c;
    input REF_CLK_c_enable_1606;
    input n31476;
    input n19_adj_1;
    output n5_adj_2;
    input n16_adj_3;
    output n17_adj_4;
    input n16_adj_5;
    output n22;
    input n16_adj_6;
    output n22_adj_7;
    input n8;
    output n2;
    input n16_adj_8;
    output n22_adj_9;
    input n16_adj_10;
    output n22_adj_11;
    input n8_adj_12;
    output n2_adj_13;
    input n41344;
    input n19_adj_14;
    output n26;
    input n359;
    output n392;
    input n16_adj_15;
    output n17_adj_16;
    input n16_adj_17;
    output n17_adj_18;
    input n17_adj_19;
    output n5_adj_20;
    input n13;
    output n14;
    input REF_CLK_c_enable_1550;
    input n41328;
    output inst1_FIFOfifo_rst;
    input REF_CLK_c_enable_1581;
    output write_ack;
    input write_ack_N_4649;
    input inst3_Empty;
    output fiford_reg;
    input fiford;
    input n40677;
    input \SHAREDBUS_ADR_I[23] ;
    input \SHAREDBUS_ADR_I[18] ;
    output n32798;
    input [31:0]inst3_Q;
    input n41347;
    output n31779;
    input n41329;
    input n41330;
    input n41331;
    input n41332;
    input n41333;
    input n41334;
    input n41335;
    input REF_CLK_c_enable_1558;
    input \SHAREDBUS_DAT_I[8] ;
    input \SHAREDBUS_DAT_I[9] ;
    input \SHAREDBUS_DAT_I[10] ;
    input \SHAREDBUS_DAT_I[11] ;
    input \SHAREDBUS_DAT_I[12] ;
    input \SHAREDBUS_DAT_I[13] ;
    input \SHAREDBUS_DAT_I[14] ;
    input \SHAREDBUS_DAT_I[15] ;
    input REF_CLK_c_enable_1566;
    input n41336;
    input n41337;
    input n41338;
    input n41339;
    input n41340;
    input n41341;
    input n41342;
    input n41343;
    input REF_CLK_c_enable_1574;
    input \SHAREDBUS_DAT_I[24] ;
    input \SHAREDBUS_DAT_I[25] ;
    input \SHAREDBUS_DAT_I[26] ;
    input \SHAREDBUS_DAT_I[27] ;
    input \SHAREDBUS_DAT_I[28] ;
    input \SHAREDBUS_DAT_I[29] ;
    input \SHAREDBUS_DAT_I[30] ;
    input \SHAREDBUS_DAT_I[31] ;
    output \reg_12[2] ;
    output \reg_12[3] ;
    output \reg_12[4] ;
    output \reg_12[6] ;
    output \reg_12[7] ;
    input REF_CLK_c_enable_1589;
    output \reg_12[9] ;
    output \reg_12[11] ;
    output \reg_12[12] ;
    output \reg_12[13] ;
    output \reg_12[14] ;
    output \reg_12[15] ;
    input REF_CLK_c_enable_1597;
    output \reg_12[17] ;
    output \reg_12[18] ;
    output \reg_12[21] ;
    output \reg_12[22] ;
    output \reg_12[24] ;
    input REF_CLK_c_enable_1605;
    output \reg_12[25] ;
    output \reg_12[28] ;
    output \reg_12[29] ;
    input inst3_Full;
    input n41193;
    input n2_adj_21;
    input n37903;
    input n2_adj_22;
    input n37905;
    input n2_adj_23;
    output n4893;
    input n2_adj_24;
    input n2_adj_25;
    input n2_adj_26;
    input n2_adj_27;
    input n37904;
    input n2_adj_28;
    input n2_adj_29;
    output n4883;
    input n2_adj_30;
    input n2_adj_31;
    output n4880;
    input n2_adj_32;
    input n2_adj_33;
    input n37906;
    input n2_adj_34;
    output n4875;
    input n2_adj_35;
    output n4873;
    input n2_adj_36;
    input n41275;
    input REF_CLK_c_enable_424;
    input n41310;
    input n30762;
    output n30241;
    output n41180;
    output n41181;
    output \FIFOwb_DAT_O[12] ;
    input n2_adj_37;
    input n2_adj_38;
    output n4868;
    input [0:0]n954;
    input [0:0]n953;
    input n41301;
    output n32366;
    input n41262;
    input n41278;
    output n35136;
    output n33088;
    input n41304;
    output n34742;
    output n41226;
    input n41255;
    input n41323;
    output n5_adj_39;
    input spiSPI_ACK_O;
    output n35042;
    input n352;
    output n385;
    input n19_adj_40;
    output n26_adj_41;
    input n19_adj_42;
    output n25;
    input n19_adj_43;
    output n25_adj_44;
    input n355;
    output n388;
    input n19_adj_45;
    output n5_adj_46;
    input n19_adj_47;
    output n25_adj_48;
    input n17_adj_49;
    output n22_adj_50;
    input n8_adj_51;
    output n2_adj_52;
    input n19_adj_53;
    output n25_adj_54;
    input n19_adj_55;
    output n25_adj_56;
    input n360;
    output n393;
    input n31183;
    input n23;
    output n31;
    input n19_adj_57;
    output n5_adj_58;
    input n8_adj_59;
    output n2_adj_60;
    input n19_adj_61;
    output n25_adj_62;
    input n19_adj_63;
    output n5_adj_64;
    output n33846;
    output \FIFOwb_DAT_O[0] ;
    input n41210;
    input n33864;
    input n19_adj_65;
    output n41258;
    output n30949;
    input \SHAREDBUS_ADR_I[30] ;
    output n41272;
    input n41265;
    output n30951;
    output n30948;
    output n30944;
    input \SHAREDBUS_ADR_I[20] ;
    input \SHAREDBUS_ADR_I[26] ;
    input \SHAREDBUS_ADR_I[27] ;
    input \SHAREDBUS_ADR_I[22] ;
    output n35844;
    output n35866;
    output n41274;
    input \SHAREDBUS_ADR_I[5] ;
    input n41346;
    output n41225;
    output n35633;
    output n35736;
    output n41277;
    input n41289;
    output n32814;
    output n35796;
    output \FIFOwb_DAT_O[18] ;
    output \FIFOwb_DAT_O[25] ;
    input n37954;
    output \FIFOwb_DAT_O[31] ;
    input n37956;
    output \FIFOwb_DAT_O[30] ;
    input n37955;
    output \FIFOwb_DAT_O[27] ;
    output \FIFOwb_DAT_O[26] ;
    output \FIFOwb_DAT_O[23] ;
    output \FIFOwb_DAT_O[20] ;
    output \FIFOwb_DAT_O[19] ;
    output \FIFOwb_DAT_O[16] ;
    output \FIFOwb_DAT_O[10] ;
    output \FIFOwb_DAT_O[8] ;
    output \FIFOwb_DAT_O[5] ;
    output \FIFOwb_DAT_O[1] ;
    output \FIFOwb_DAT_O[21] ;
    output \FIFOwb_DAT_O[28] ;
    output \FIFOwb_DAT_O[15] ;
    output \FIFOwb_DAT_O[13] ;
    output \FIFOwb_DAT_O[11] ;
    output \FIFOwb_DAT_O[9] ;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    
    wire n32820, n32812, n41261;
    wire [31:0]status_reg;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(111[15:25])
    wire [31:0]reg_12;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(106[15:21])
    
    wire n36170, n36112, n36113, n36114;
    wire [7:0]FIFOout_pins;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/platform1_vhd.vhd(16[3:15])
    
    wire n40678, n40679;
    wire [31:0]reg_00;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(103[15:21])
    
    wire n1, n1_adj_5839, n1_adj_5840, n1_adj_5841, n1_adj_5842, n1_adj_5843, 
        n1_adj_5844, n1_adj_5845, n1_adj_5846, n1_adj_5847, n1_adj_5848, 
        n1_adj_5849, n1_adj_5850, n1_adj_5851, n1_adj_5852, n1_adj_5853, 
        n1_adj_5854, n1_adj_5855, n36169, n1_adj_5856;
    wire [31:0]n4865;
    
    wire n1_adj_5857, n1_adj_5858, n1_adj_5859, n1_adj_5860, n1_adj_5861, 
        n1_adj_5862, n1_adj_5863, n1_adj_5864, n1_adj_5865, n1_adj_5866, 
        n36171, n33878, n33870, n41290, n33858, n33802, n33720, 
        n33788, n33784, n33894;
    
    LUT4 i1_4_lut (.A(n32828), .B(n41246), .C(n34372), .D(n32820), .Z(n5223)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 i1_4_lut_adj_202 (.A(n15), .B(n32812), .C(n41261), .D(n41303), 
         .Z(n32820)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_202.init = 16'hfffe;
    LUT4 i1_4_lut_adj_203 (.A(\SHAREDBUS_ADR_I[25] ), .B(\SHAREDBUS_ADR_I[24] ), 
         .C(\SHAREDBUS_ADR_I[29] ), .D(\SHAREDBUS_ADR_I[16] ), .Z(n32812)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_203.init = 16'hfffe;
    LUT4 i30998_3_lut (.A(status_reg[1]), .B(reg_12[1]), .C(n41345), .Z(n36170)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30998_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n16), 
         .Z(n17)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_204 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n19), 
         .Z(n5)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_204.init = 16'hd0d0;
    FD1S3DX read_ack_153 (.D(n31476), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(read_ack)) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(153[12] 160[10])
    defparam read_ack_153.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_205 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n19_adj_1), 
         .Z(n5_adj_2)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_205.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_206 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n16_adj_3), 
         .Z(n17_adj_4)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_206.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_207 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n16_adj_5), 
         .Z(n22)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_207.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_208 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n16_adj_6), 
         .Z(n22_adj_7)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_208.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_209 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n8), 
         .Z(n2)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_209.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_210 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n16_adj_8), 
         .Z(n22_adj_9)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_210.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_211 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n16_adj_10), 
         .Z(n22_adj_11)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_211.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_212 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n8_adj_12), 
         .Z(n2_adj_13)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_212.init = 16'hd0d0;
    PFUMX i30942 (.BLUT(n36112), .ALUT(n36113), .C0(n41344), .Z(n36114));
    LUT4 i1_2_lut_3_lut_adj_213 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n19_adj_14), 
         .Z(n26)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_213.init = 16'hd0d0;
    LUT4 i14845_2_lut_3_lut (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n359), 
         .Z(n392)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i14845_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_214 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n16_adj_15), 
         .Z(n17_adj_16)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_214.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_215 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n16_adj_17), 
         .Z(n17_adj_18)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_215.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_216 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n17_adj_19), 
         .Z(n5_adj_20)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_216.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_217 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n13), 
         .Z(n14)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_217.init = 16'he0e0;
    FD1P3DX reg_00__i1 (.D(n41328), .SP(REF_CLK_c_enable_1550), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(FIFOout_pins[0])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i1.GSR = "ENABLED";
    FD1P3DX reg_12__i0 (.D(n41328), .SP(REF_CLK_c_enable_1581), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(inst1_FIFOfifo_rst)) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i0.GSR = "ENABLED";
    FD1S3DX write_ack_154 (.D(write_ack_N_4649), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(write_ack)) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(178[12] 186[10])
    defparam write_ack_154.GSR = "ENABLED";
    FD1S3DX status_reg_i1 (.D(inst3_Empty), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(status_reg[0])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(195[12] 199[10])
    defparam status_reg_i1.GSR = "ENABLED";
    FD1S3DX fiford_reg_156 (.D(fiford), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(fiford_reg)) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(210[12] 212[10])
    defparam fiford_reg_156.GSR = "ENABLED";
    PFUMX i34154 (.BLUT(n40678), .ALUT(n40677), .C0(n41344), .Z(n40679));
    LUT4 i1_2_lut (.A(\SHAREDBUS_ADR_I[23] ), .B(\SHAREDBUS_ADR_I[18] ), 
         .Z(n32798)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 mux_1642_Mux_29_i1_3_lut (.A(reg_00[29]), .B(inst3_Q[29]), .C(n41345), 
         .Z(n1)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_29_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_28_i1_3_lut (.A(reg_00[28]), .B(inst3_Q[28]), .C(n41345), 
         .Z(n1_adj_5839)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_28_i1_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut (.A(n41344), .B(n41345), .C(n41347), .Z(n31779)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_3_lut.init = 16'hfbfb;
    LUT4 mux_1642_Mux_25_i1_3_lut (.A(reg_00[25]), .B(inst3_Q[25]), .C(n41345), 
         .Z(n1_adj_5840)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_25_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_24_i1_3_lut (.A(reg_00[24]), .B(inst3_Q[24]), .C(n41345), 
         .Z(n1_adj_5841)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_24_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_22_i1_3_lut (.A(reg_00[22]), .B(inst3_Q[22]), .C(n41345), 
         .Z(n1_adj_5842)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_22_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_21_i1_3_lut (.A(reg_00[21]), .B(inst3_Q[21]), .C(n41345), 
         .Z(n1_adj_5843)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_21_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_18_i1_3_lut (.A(reg_00[18]), .B(inst3_Q[18]), .C(n41345), 
         .Z(n1_adj_5844)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_18_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_17_i1_3_lut (.A(reg_00[17]), .B(inst3_Q[17]), .C(n41345), 
         .Z(n1_adj_5845)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_17_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_15_i1_3_lut (.A(reg_00[15]), .B(inst3_Q[15]), .C(n41345), 
         .Z(n1_adj_5846)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_15_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_14_i1_3_lut (.A(reg_00[14]), .B(inst3_Q[14]), .C(n41345), 
         .Z(n1_adj_5847)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_14_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_13_i1_3_lut (.A(reg_00[13]), .B(inst3_Q[13]), .C(n41345), 
         .Z(n1_adj_5848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_13_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_11_i1_3_lut (.A(reg_00[11]), .B(inst3_Q[11]), .C(n41345), 
         .Z(n1_adj_5849)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_11_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_9_i1_3_lut (.A(reg_00[9]), .B(inst3_Q[9]), .C(n41345), 
         .Z(n1_adj_5850)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_9_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_7_i1_3_lut (.A(FIFOout_pins[7]), .B(inst3_Q[7]), .C(n41345), 
         .Z(n1_adj_5851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_7_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_6_i1_3_lut (.A(FIFOout_pins[6]), .B(inst3_Q[6]), .C(n41345), 
         .Z(n1_adj_5852)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_6_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_4_i1_3_lut (.A(FIFOout_pins[4]), .B(inst3_Q[4]), .C(n41345), 
         .Z(n1_adj_5853)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_4_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_3_i1_3_lut (.A(FIFOout_pins[3]), .B(inst3_Q[3]), .C(n41345), 
         .Z(n1_adj_5854)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_3_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_2_i1_3_lut (.A(FIFOout_pins[2]), .B(inst3_Q[2]), .C(n41345), 
         .Z(n1_adj_5855)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_2_i1_3_lut.init = 16'hcaca;
    FD1P3DX reg_00__i2 (.D(n41329), .SP(REF_CLK_c_enable_1550), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(FIFOout_pins[1])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i2.GSR = "ENABLED";
    FD1P3DX reg_00__i3 (.D(n41330), .SP(REF_CLK_c_enable_1550), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(FIFOout_pins[2])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i3.GSR = "ENABLED";
    FD1P3DX reg_00__i4 (.D(n41331), .SP(REF_CLK_c_enable_1550), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(FIFOout_pins[3])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i4.GSR = "ENABLED";
    FD1P3DX reg_00__i5 (.D(n41332), .SP(REF_CLK_c_enable_1550), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(FIFOout_pins[4])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i5.GSR = "ENABLED";
    FD1P3DX reg_00__i6 (.D(n41333), .SP(REF_CLK_c_enable_1550), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(FIFOout_pins[5])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i6.GSR = "ENABLED";
    FD1P3DX reg_00__i7 (.D(n41334), .SP(REF_CLK_c_enable_1550), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(FIFOout_pins[6])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i7.GSR = "ENABLED";
    FD1P3DX reg_00__i8 (.D(n41335), .SP(REF_CLK_c_enable_1550), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(FIFOout_pins[7])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i8.GSR = "ENABLED";
    FD1P3DX reg_00__i9 (.D(\SHAREDBUS_DAT_I[8] ), .SP(REF_CLK_c_enable_1558), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[8])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i9.GSR = "ENABLED";
    FD1P3DX reg_00__i10 (.D(\SHAREDBUS_DAT_I[9] ), .SP(REF_CLK_c_enable_1558), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[9])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i10.GSR = "ENABLED";
    FD1P3DX reg_00__i11 (.D(\SHAREDBUS_DAT_I[10] ), .SP(REF_CLK_c_enable_1558), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[10])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i11.GSR = "ENABLED";
    FD1P3DX reg_00__i12 (.D(\SHAREDBUS_DAT_I[11] ), .SP(REF_CLK_c_enable_1558), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[11])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i12.GSR = "ENABLED";
    FD1P3DX reg_00__i13 (.D(\SHAREDBUS_DAT_I[12] ), .SP(REF_CLK_c_enable_1558), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[12])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i13.GSR = "ENABLED";
    FD1P3DX reg_00__i14 (.D(\SHAREDBUS_DAT_I[13] ), .SP(REF_CLK_c_enable_1558), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[13])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i14.GSR = "ENABLED";
    FD1P3DX reg_00__i15 (.D(\SHAREDBUS_DAT_I[14] ), .SP(REF_CLK_c_enable_1558), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[14])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i15.GSR = "ENABLED";
    FD1P3DX reg_00__i16 (.D(\SHAREDBUS_DAT_I[15] ), .SP(REF_CLK_c_enable_1558), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[15])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i16.GSR = "ENABLED";
    FD1P3DX reg_00__i17 (.D(n41336), .SP(REF_CLK_c_enable_1566), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_00[16])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i17.GSR = "ENABLED";
    FD1P3DX reg_00__i18 (.D(n41337), .SP(REF_CLK_c_enable_1566), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_00[17])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i18.GSR = "ENABLED";
    FD1P3DX reg_00__i19 (.D(n41338), .SP(REF_CLK_c_enable_1566), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_00[18])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i19.GSR = "ENABLED";
    FD1P3DX reg_00__i20 (.D(n41339), .SP(REF_CLK_c_enable_1566), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_00[19])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i20.GSR = "ENABLED";
    FD1P3DX reg_00__i21 (.D(n41340), .SP(REF_CLK_c_enable_1566), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_00[20])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i21.GSR = "ENABLED";
    FD1P3DX reg_00__i22 (.D(n41341), .SP(REF_CLK_c_enable_1566), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_00[21])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i22.GSR = "ENABLED";
    FD1P3DX reg_00__i23 (.D(n41342), .SP(REF_CLK_c_enable_1566), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_00[22])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i23.GSR = "ENABLED";
    FD1P3DX reg_00__i24 (.D(n41343), .SP(REF_CLK_c_enable_1566), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_00[23])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i24.GSR = "ENABLED";
    FD1P3DX reg_00__i25 (.D(\SHAREDBUS_DAT_I[24] ), .SP(REF_CLK_c_enable_1574), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[24])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i25.GSR = "ENABLED";
    FD1P3DX reg_00__i26 (.D(\SHAREDBUS_DAT_I[25] ), .SP(REF_CLK_c_enable_1574), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[25])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i26.GSR = "ENABLED";
    FD1P3DX reg_00__i27 (.D(\SHAREDBUS_DAT_I[26] ), .SP(REF_CLK_c_enable_1574), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[26])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i27.GSR = "ENABLED";
    FD1P3DX reg_00__i28 (.D(\SHAREDBUS_DAT_I[27] ), .SP(REF_CLK_c_enable_1574), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[27])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i28.GSR = "ENABLED";
    FD1P3DX reg_00__i29 (.D(\SHAREDBUS_DAT_I[28] ), .SP(REF_CLK_c_enable_1574), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[28])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i29.GSR = "ENABLED";
    FD1P3DX reg_00__i30 (.D(\SHAREDBUS_DAT_I[29] ), .SP(REF_CLK_c_enable_1574), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[29])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i30.GSR = "ENABLED";
    FD1P3DX reg_00__i31 (.D(\SHAREDBUS_DAT_I[30] ), .SP(REF_CLK_c_enable_1574), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[30])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i31.GSR = "ENABLED";
    FD1P3DX reg_00__i32 (.D(\SHAREDBUS_DAT_I[31] ), .SP(REF_CLK_c_enable_1574), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_00[31])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(221[12] 237[10])
    defparam reg_00__i32.GSR = "ENABLED";
    FD1P3DX reg_12__i1 (.D(n41329), .SP(REF_CLK_c_enable_1581), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_12[1])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i1.GSR = "ENABLED";
    FD1P3DX reg_12__i2 (.D(n41330), .SP(REF_CLK_c_enable_1581), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_12[2] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i2.GSR = "ENABLED";
    FD1P3DX reg_12__i3 (.D(n41331), .SP(REF_CLK_c_enable_1581), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_12[3] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i3.GSR = "ENABLED";
    FD1P3DX reg_12__i4 (.D(n41332), .SP(REF_CLK_c_enable_1581), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_12[4] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i4.GSR = "ENABLED";
    FD1P3DX reg_12__i5 (.D(n41333), .SP(REF_CLK_c_enable_1581), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_12[5])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i5.GSR = "ENABLED";
    FD1P3DX reg_12__i6 (.D(n41334), .SP(REF_CLK_c_enable_1581), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_12[6] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i6.GSR = "ENABLED";
    FD1P3DX reg_12__i7 (.D(n41335), .SP(REF_CLK_c_enable_1581), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_12[7] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i7.GSR = "ENABLED";
    FD1P3DX reg_12__i8 (.D(\SHAREDBUS_DAT_I[8] ), .SP(REF_CLK_c_enable_1589), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_12[8])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i8.GSR = "ENABLED";
    FD1P3DX reg_12__i9 (.D(\SHAREDBUS_DAT_I[9] ), .SP(REF_CLK_c_enable_1589), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_12[9] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i9.GSR = "ENABLED";
    FD1P3DX reg_12__i10 (.D(\SHAREDBUS_DAT_I[10] ), .SP(REF_CLK_c_enable_1589), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_12[10])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i10.GSR = "ENABLED";
    FD1P3DX reg_12__i11 (.D(\SHAREDBUS_DAT_I[11] ), .SP(REF_CLK_c_enable_1589), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_12[11] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i11.GSR = "ENABLED";
    FD1P3DX reg_12__i12 (.D(\SHAREDBUS_DAT_I[12] ), .SP(REF_CLK_c_enable_1589), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_12[12] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i12.GSR = "ENABLED";
    FD1P3DX reg_12__i13 (.D(\SHAREDBUS_DAT_I[13] ), .SP(REF_CLK_c_enable_1589), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_12[13] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i13.GSR = "ENABLED";
    FD1P3DX reg_12__i14 (.D(\SHAREDBUS_DAT_I[14] ), .SP(REF_CLK_c_enable_1589), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_12[14] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i14.GSR = "ENABLED";
    FD1P3DX reg_12__i15 (.D(\SHAREDBUS_DAT_I[15] ), .SP(REF_CLK_c_enable_1589), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_12[15] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i15.GSR = "ENABLED";
    FD1P3DX reg_12__i16 (.D(n41336), .SP(REF_CLK_c_enable_1597), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_12[16])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i16.GSR = "ENABLED";
    FD1P3DX reg_12__i17 (.D(n41337), .SP(REF_CLK_c_enable_1597), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_12[17] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i17.GSR = "ENABLED";
    FD1P3DX reg_12__i18 (.D(n41338), .SP(REF_CLK_c_enable_1597), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_12[18] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i18.GSR = "ENABLED";
    FD1P3DX reg_12__i19 (.D(n41339), .SP(REF_CLK_c_enable_1597), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_12[19])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i19.GSR = "ENABLED";
    FD1P3DX reg_12__i20 (.D(n41340), .SP(REF_CLK_c_enable_1597), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_12[20])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i20.GSR = "ENABLED";
    FD1P3DX reg_12__i21 (.D(n41341), .SP(REF_CLK_c_enable_1597), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_12[21] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i21.GSR = "ENABLED";
    FD1P3DX reg_12__i22 (.D(n41342), .SP(REF_CLK_c_enable_1597), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(\reg_12[22] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i22.GSR = "ENABLED";
    FD1P3DX reg_12__i23 (.D(n41343), .SP(REF_CLK_c_enable_1597), .CK(REF_CLK_c), 
            .CD(REF_CLK_c_enable_1606), .Q(reg_12[23])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i23.GSR = "ENABLED";
    FD1P3DX reg_12__i24 (.D(\SHAREDBUS_DAT_I[24] ), .SP(REF_CLK_c_enable_1605), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_12[24] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i24.GSR = "ENABLED";
    FD1P3DX reg_12__i25 (.D(\SHAREDBUS_DAT_I[25] ), .SP(REF_CLK_c_enable_1605), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_12[25] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i25.GSR = "ENABLED";
    FD1P3DX reg_12__i26 (.D(\SHAREDBUS_DAT_I[26] ), .SP(REF_CLK_c_enable_1605), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_12[26])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i26.GSR = "ENABLED";
    FD1P3DX reg_12__i27 (.D(\SHAREDBUS_DAT_I[27] ), .SP(REF_CLK_c_enable_1605), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_12[27])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i27.GSR = "ENABLED";
    FD1P3DX reg_12__i28 (.D(\SHAREDBUS_DAT_I[28] ), .SP(REF_CLK_c_enable_1605), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_12[28] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i28.GSR = "ENABLED";
    FD1P3DX reg_12__i29 (.D(\SHAREDBUS_DAT_I[29] ), .SP(REF_CLK_c_enable_1605), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(\reg_12[29] )) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i29.GSR = "ENABLED";
    FD1P3DX reg_12__i30 (.D(\SHAREDBUS_DAT_I[30] ), .SP(REF_CLK_c_enable_1605), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_12[30])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i30.GSR = "ENABLED";
    FD1P3DX reg_12__i31 (.D(\SHAREDBUS_DAT_I[31] ), .SP(REF_CLK_c_enable_1605), 
            .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), .Q(reg_12[31])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(246[12] 262[10])
    defparam reg_12__i31.GSR = "ENABLED";
    FD1S3DX status_reg_i2 (.D(inst3_Full), .CK(REF_CLK_c), .CD(REF_CLK_c_enable_1606), 
            .Q(status_reg[1])) /* synthesis LSE_LINE_FILE_ID=41, LSE_LCOL=11, LSE_RCOL=34, LSE_LLINE=83, LSE_RLINE=109 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(195[12] 199[10])
    defparam status_reg_i2.GSR = "ENABLED";
    LUT4 i30997_3_lut (.A(FIFOout_pins[1]), .B(inst3_Q[1]), .C(n41345), 
         .Z(n36169)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30997_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_5_i1_3_lut (.A(FIFOout_pins[5]), .B(inst3_Q[5]), .C(n41345), 
         .Z(n1_adj_5856)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_5_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_8_i3_4_lut (.A(reg_12[8]), .B(n41193), .C(n5223), 
         .D(n41345), .Z(n4865[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_8_i3_4_lut.init = 16'hcac0;
    LUT4 mux_1642_Mux_8_i1_3_lut (.A(reg_00[8]), .B(inst3_Q[8]), .C(n41345), 
         .Z(n1_adj_5857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_8_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_10_i1_3_lut (.A(reg_00[10]), .B(inst3_Q[10]), .C(n41345), 
         .Z(n1_adj_5858)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_10_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_16_i1_3_lut (.A(reg_00[16]), .B(inst3_Q[16]), .C(n41345), 
         .Z(n1_adj_5859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_16_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_19_i1_3_lut (.A(reg_00[19]), .B(inst3_Q[19]), .C(n41345), 
         .Z(n1_adj_5860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_19_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_20_i3_4_lut (.A(reg_12[20]), .B(n41193), .C(n5223), 
         .D(n41345), .Z(n4865[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_20_i3_4_lut.init = 16'hcac0;
    LUT4 mux_1642_Mux_20_i1_3_lut (.A(reg_00[20]), .B(inst3_Q[20]), .C(n41345), 
         .Z(n1_adj_5861)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_20_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_23_i1_3_lut (.A(reg_00[23]), .B(inst3_Q[23]), .C(n41345), 
         .Z(n1_adj_5862)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_23_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_26_i1_3_lut (.A(reg_00[26]), .B(inst3_Q[26]), .C(n41345), 
         .Z(n1_adj_5863)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_26_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_27_i1_3_lut (.A(reg_00[27]), .B(inst3_Q[27]), .C(n41345), 
         .Z(n1_adj_5864)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_27_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_30_i1_3_lut (.A(reg_00[30]), .B(inst3_Q[30]), .C(n41345), 
         .Z(n1_adj_5865)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_30_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1642_Mux_31_i1_3_lut (.A(reg_00[31]), .B(inst3_Q[31]), .C(n41345), 
         .Z(n1_adj_5866)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(165[25] 170[37])
    defparam mux_1642_Mux_31_i1_3_lut.init = 16'hcaca;
    PFUMX mux_1642_Mux_2_i3 (.BLUT(n1_adj_5855), .ALUT(n2_adj_21), .C0(n37903), 
          .Z(n4865[2]));
    PFUMX mux_1642_Mux_3_i3 (.BLUT(n1_adj_5854), .ALUT(n2_adj_22), .C0(n37905), 
          .Z(n4865[3]));
    PFUMX mux_1642_Mux_4_i3 (.BLUT(n1_adj_5853), .ALUT(n2_adj_23), .C0(n37905), 
          .Z(n4893));
    PFUMX mux_1642_Mux_6_i3 (.BLUT(n1_adj_5852), .ALUT(n2_adj_24), .C0(n37905), 
          .Z(n4865[6]));
    PFUMX mux_1642_Mux_7_i3 (.BLUT(n1_adj_5851), .ALUT(n2_adj_25), .C0(n37905), 
          .Z(n4865[7]));
    PFUMX mux_1642_Mux_9_i3 (.BLUT(n1_adj_5850), .ALUT(n2_adj_26), .C0(n37903), 
          .Z(n4865[9]));
    PFUMX mux_1642_Mux_11_i3 (.BLUT(n1_adj_5849), .ALUT(n2_adj_27), .C0(n37904), 
          .Z(n4865[11]));
    PFUMX mux_1642_Mux_13_i3 (.BLUT(n1_adj_5848), .ALUT(n2_adj_28), .C0(n37903), 
          .Z(n4865[13]));
    PFUMX mux_1642_Mux_14_i3 (.BLUT(n1_adj_5847), .ALUT(n2_adj_29), .C0(n37904), 
          .Z(n4883));
    PFUMX mux_1642_Mux_15_i3 (.BLUT(n1_adj_5846), .ALUT(n2_adj_30), .C0(n37903), 
          .Z(n4865[15]));
    PFUMX mux_1642_Mux_17_i3 (.BLUT(n1_adj_5845), .ALUT(n2_adj_31), .C0(n37904), 
          .Z(n4880));
    PFUMX mux_1642_Mux_18_i3 (.BLUT(n1_adj_5844), .ALUT(n2_adj_32), .C0(n37904), 
          .Z(n4865[18]));
    PFUMX mux_1642_Mux_21_i3 (.BLUT(n1_adj_5843), .ALUT(n2_adj_33), .C0(n37906), 
          .Z(n4865[21]));
    PFUMX mux_1642_Mux_22_i3 (.BLUT(n1_adj_5842), .ALUT(n2_adj_34), .C0(n37906), 
          .Z(n4875));
    PFUMX mux_1642_Mux_24_i3 (.BLUT(n1_adj_5841), .ALUT(n2_adj_35), .C0(n37906), 
          .Z(n4873));
    PFUMX mux_1642_Mux_25_i3 (.BLUT(n1_adj_5840), .ALUT(n2_adj_36), .C0(n37906), 
          .Z(n4865[25]));
    LUT4 i25224_2_lut_4_lut (.A(n41275), .B(REF_CLK_c_enable_424), .C(n41310), 
         .D(n30762), .Z(n30241)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i25224_2_lut_4_lut.init = 16'h00fb;
    LUT4 i33275_2_lut_rep_775_4_lut (.A(n41275), .B(REF_CLK_c_enable_424), 
         .C(n41310), .D(\SHAREDBUS_ADR_I[7] ), .Z(n41180)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i33275_2_lut_rep_775_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_rep_776_4_lut (.A(n41275), .B(REF_CLK_c_enable_424), .C(n41310), 
         .D(\SHAREDBUS_ADR_I[7] ), .Z(n41181)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_rep_776_4_lut.init = 16'hfffb;
    LUT4 i30999_3_lut_3_lut (.A(n41193), .B(n5223), .C(n36170), .Z(n36171)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(169[25] 170[37])
    defparam i30999_3_lut_3_lut.init = 16'h7474;
    LUT4 n40679_bdd_3_lut_3_lut (.A(n41193), .B(n5223), .C(n40679), .Z(\FIFOwb_DAT_O[12] )) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(169[25] 170[37])
    defparam n40679_bdd_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_1642_Mux_31_i3_4_lut_4_lut (.A(n41193), .B(n41345), .C(n5223), 
         .D(reg_12[31]), .Z(n4865[31])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(169[25] 170[37])
    defparam mux_1642_Mux_31_i3_4_lut_4_lut.init = 16'h5c50;
    LUT4 mux_1642_Mux_30_i3_4_lut_4_lut (.A(n41193), .B(n41345), .C(n5223), 
         .D(reg_12[30]), .Z(n4865[30])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(169[25] 170[37])
    defparam mux_1642_Mux_30_i3_4_lut_4_lut.init = 16'h5c50;
    LUT4 mux_1642_Mux_26_i3_4_lut_4_lut (.A(n41193), .B(n41345), .C(n5223), 
         .D(reg_12[26]), .Z(n4865[26])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(169[25] 170[37])
    defparam mux_1642_Mux_26_i3_4_lut_4_lut.init = 16'h5c50;
    LUT4 mux_1642_Mux_23_i3_4_lut_4_lut (.A(n41193), .B(n41345), .C(n5223), 
         .D(reg_12[23]), .Z(n4865[23])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(169[25] 170[37])
    defparam mux_1642_Mux_23_i3_4_lut_4_lut.init = 16'h5c50;
    LUT4 mux_1642_Mux_19_i3_4_lut_4_lut (.A(n41193), .B(n41345), .C(n5223), 
         .D(reg_12[19]), .Z(n4865[19])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(169[25] 170[37])
    defparam mux_1642_Mux_19_i3_4_lut_4_lut.init = 16'h5c50;
    LUT4 mux_1642_Mux_16_i3_4_lut_4_lut (.A(n41193), .B(n41345), .C(n5223), 
         .D(reg_12[16]), .Z(n4865[16])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(169[25] 170[37])
    defparam mux_1642_Mux_16_i3_4_lut_4_lut.init = 16'h5c50;
    LUT4 mux_1642_Mux_10_i3_4_lut_4_lut (.A(n41193), .B(n41345), .C(n5223), 
         .D(reg_12[10]), .Z(n4865[10])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(169[25] 170[37])
    defparam mux_1642_Mux_10_i3_4_lut_4_lut.init = 16'h5c50;
    LUT4 mux_1642_Mux_5_i3_4_lut_4_lut (.A(n41193), .B(n41345), .C(n5223), 
         .D(reg_12[5]), .Z(n4865[5])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(169[25] 170[37])
    defparam mux_1642_Mux_5_i3_4_lut_4_lut.init = 16'h5c50;
    LUT4 mux_1642_Mux_27_i3_4_lut_4_lut (.A(n41193), .B(n41345), .C(n5223), 
         .D(reg_12[27]), .Z(n4865[27])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(169[25] 170[37])
    defparam mux_1642_Mux_27_i3_4_lut_4_lut.init = 16'h5c50;
    PFUMX mux_1642_Mux_28_i3 (.BLUT(n1_adj_5839), .ALUT(n2_adj_37), .C0(n41344), 
          .Z(n4865[28]));
    PFUMX mux_1642_Mux_29_i3 (.BLUT(n1), .ALUT(n2_adj_38), .C0(n41344), 
          .Z(n4868));
    LUT4 i1_2_lut_rep_841 (.A(n954[0]), .B(n953[0]), .Z(n41246)) /* synthesis lut_function=(A (B)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(137[25:61])
    defparam i1_2_lut_rep_841.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_218 (.A(n954[0]), .B(n953[0]), .C(n41301), 
         .Z(n32366)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(137[25:61])
    defparam i1_2_lut_3_lut_adj_218.init = 16'h8080;
    LUT4 i1_3_lut_4_lut (.A(n954[0]), .B(n953[0]), .C(n41262), .D(n41278), 
         .Z(n35136)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(137[25:61])
    defparam i1_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_3_lut_4_lut_adj_219 (.A(n954[0]), .B(n953[0]), .C(n41262), 
         .D(n41303), .Z(n33088)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(137[25:61])
    defparam i1_3_lut_4_lut_adj_219.init = 16'h0080;
    LUT4 i1_3_lut_4_lut_adj_220 (.A(n954[0]), .B(n953[0]), .C(n41310), 
         .D(n41304), .Z(n34742)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(137[25:61])
    defparam i1_3_lut_4_lut_adj_220.init = 16'h0080;
    LUT4 i1_3_lut_rep_821_4_lut (.A(n954[0]), .B(n953[0]), .C(n41303), 
         .D(n41347), .Z(n41226)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(137[25:61])
    defparam i1_3_lut_rep_821_4_lut.init = 16'h0008;
    LUT4 i1_3_lut_4_lut_adj_221 (.A(n954[0]), .B(n953[0]), .C(n41255), 
         .D(n41323), .Z(n5_adj_39)) /* synthesis lut_function=(A (B (C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(137[25:61])
    defparam i1_3_lut_4_lut_adj_221.init = 16'h8088;
    LUT4 i1_3_lut_4_lut_adj_222 (.A(n954[0]), .B(n953[0]), .C(spiSPI_ACK_O), 
         .D(n41310), .Z(n35042)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(137[25:61])
    defparam i1_3_lut_4_lut_adj_222.init = 16'h0800;
    LUT4 i14847_2_lut_3_lut (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n352), 
         .Z(n385)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i14847_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_223 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n19_adj_40), 
         .Z(n26_adj_41)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_223.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_224 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n19_adj_42), 
         .Z(n25)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_224.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_225 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n19_adj_43), 
         .Z(n25_adj_44)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_225.init = 16'hd0d0;
    LUT4 i14846_2_lut_3_lut (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n355), 
         .Z(n388)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i14846_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_226 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n19_adj_45), 
         .Z(n5_adj_46)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_226.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_227 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n19_adj_47), 
         .Z(n25_adj_48)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_227.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_228 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n17_adj_49), 
         .Z(n22_adj_50)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_228.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_229 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n8_adj_51), 
         .Z(n2_adj_52)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_229.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_230 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n19_adj_53), 
         .Z(n25_adj_54)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_230.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_231 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n19_adj_55), 
         .Z(n25_adj_56)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_231.init = 16'hd0d0;
    LUT4 i14500_2_lut_3_lut (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n360), 
         .Z(n393)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i14500_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i32942_3_lut_4_lut (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n31183), 
         .D(n23), .Z(n31)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i32942_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_3_lut_adj_232 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n19_adj_57), 
         .Z(n5_adj_58)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_232.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_233 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n8_adj_59), 
         .Z(n2_adj_60)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_233.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_234 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n19_adj_61), 
         .Z(n25_adj_62)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_234.init = 16'hd0d0;
    LUT4 i1_2_lut_3_lut_adj_235 (.A(\SHAREDBUS_ADR_I[7] ), .B(n41186), .C(n19_adj_63), 
         .Z(n5_adj_64)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_adj_235.init = 16'hd0d0;
    LUT4 i1_2_lut_adj_236 (.A(\SHAREDBUS_ADR_I[18] ), .B(\SHAREDBUS_ADR_I[25] ), 
         .Z(n33846)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_236.init = 16'heeee;
    LUT4 i1_4_lut_adj_237 (.A(n33878), .B(n41246), .C(n34372), .D(n33870), 
         .Z(\FIFOwb_DAT_O[0] )) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut_adj_237.init = 16'hfffb;
    LUT4 i1_4_lut_adj_238 (.A(n41210), .B(n33864), .C(n41310), .D(n19_adj_65), 
         .Z(n33878)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i1_4_lut_adj_238.init = 16'hffdf;
    LUT4 i1_4_lut_adj_239 (.A(n15), .B(n41290), .C(n33858), .D(n41258), 
         .Z(n33870)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_239.init = 16'hfffe;
    LUT4 i1_4_lut_adj_240 (.A(n41246), .B(n33802), .C(n4865[2]), .D(n33720), 
         .Z(n30949)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_240.init = 16'hfffd;
    LUT4 i1_4_lut_adj_241 (.A(n34372), .B(n41210), .C(n15), .D(n33788), 
         .Z(n33802)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut_adj_241.init = 16'hfffb;
    LUT4 i1_4_lut_adj_242 (.A(\SHAREDBUS_ADR_I[30] ), .B(n33784), .C(n41272), 
         .D(\SHAREDBUS_ADR_I[16] ), .Z(n33788)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_242.init = 16'hfffe;
    LUT4 i1_4_lut_adj_243 (.A(n33894), .B(n41310), .C(n19_adj_65), .D(n41265), 
         .Z(n33720)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut_adj_243.init = 16'hfffb;
    LUT4 i1_4_lut_adj_244 (.A(n41246), .B(n33802), .C(n4865[3]), .D(n33720), 
         .Z(n30951)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_244.init = 16'hfffd;
    LUT4 i1_4_lut_adj_245 (.A(n41246), .B(n33802), .C(n4865[6]), .D(n33720), 
         .Z(n30948)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_245.init = 16'hfffd;
    LUT4 i1_4_lut_adj_246 (.A(n41246), .B(n33802), .C(n4865[7]), .D(n33720), 
         .Z(n30944)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_246.init = 16'hfffd;
    LUT4 i1_2_lut_rep_853 (.A(\SHAREDBUS_ADR_I[20] ), .B(\SHAREDBUS_ADR_I[26] ), 
         .Z(n41258)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_853.init = 16'heeee;
    LUT4 i1_2_lut_rep_856 (.A(\SHAREDBUS_ADR_I[30] ), .B(\SHAREDBUS_ADR_I[27] ), 
         .Z(n41261)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_856.init = 16'heeee;
    LUT4 i30682_3_lut_4_lut (.A(\SHAREDBUS_ADR_I[30] ), .B(\SHAREDBUS_ADR_I[27] ), 
         .C(\SHAREDBUS_ADR_I[18] ), .D(\SHAREDBUS_ADR_I[22] ), .Z(n35844)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30682_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_867 (.A(\SHAREDBUS_ADR_I[25] ), .B(\SHAREDBUS_ADR_I[23] ), 
         .Z(n41272)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_867.init = 16'heeee;
    LUT4 i30704_2_lut_3_lut_4_lut (.A(\SHAREDBUS_ADR_I[25] ), .B(\SHAREDBUS_ADR_I[23] ), 
         .C(\SHAREDBUS_ADR_I[24] ), .D(\SHAREDBUS_ADR_I[18] ), .Z(n35866)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30704_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 SHAREDBUS_ADR_I_3__bdd_3_lut (.A(n41345), .B(reg_00[12]), .C(inst3_Q[12]), 
         .Z(n40678)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam SHAREDBUS_ADR_I_3__bdd_3_lut.init = 16'he4e4;
    LUT4 i1_2_lut_rep_869 (.A(\SHAREDBUS_ADR_I[30] ), .B(\SHAREDBUS_ADR_I[24] ), 
         .Z(n41274)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_869.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_247 (.A(\SHAREDBUS_ADR_I[30] ), .B(\SHAREDBUS_ADR_I[24] ), 
         .C(n36114), .D(n41347), .Z(n33858)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_247.init = 16'hfffe;
    LUT4 i1_3_lut_rep_781_4_lut (.A(\SHAREDBUS_ADR_I[5] ), .B(n41346), .C(n41310), 
         .D(REF_CLK_c_enable_424), .Z(n41186)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_3_lut_rep_781_4_lut.init = 16'hfeff;
    LUT4 i1_2_lut_rep_820_3_lut (.A(\SHAREDBUS_ADR_I[5] ), .B(n41346), .C(\SHAREDBUS_ADR_I[7] ), 
         .Z(n41225)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_rep_820_3_lut.init = 16'hfefe;
    LUT4 i30475_2_lut_3_lut_4_lut (.A(\SHAREDBUS_ADR_I[5] ), .B(n41346), 
         .C(n15), .D(\SHAREDBUS_ADR_I[7] ), .Z(n35633)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i30475_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i30577_2_lut_3_lut_4_lut (.A(\SHAREDBUS_ADR_I[5] ), .B(n41346), 
         .C(n41310), .D(\SHAREDBUS_ADR_I[7] ), .Z(n35736)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i30577_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\SHAREDBUS_ADR_I[5] ), .B(n41346), .C(n41301), 
         .D(\SHAREDBUS_ADR_I[7] ), .Z(n34372)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/platform1/soc/../components/FIFO_Comp/rtl/verilog/wb_fifo_dev.v(132[7:30])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hffef;
    LUT4 i1_2_lut_rep_872 (.A(\SHAREDBUS_ADR_I[26] ), .B(\SHAREDBUS_ADR_I[22] ), 
         .Z(n41277)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_872.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_248 (.A(\SHAREDBUS_ADR_I[26] ), .B(\SHAREDBUS_ADR_I[22] ), 
         .C(n41289), .D(n32798), .Z(n32814)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_248.init = 16'hfffe;
    LUT4 i30634_2_lut_3_lut_4_lut (.A(\SHAREDBUS_ADR_I[26] ), .B(\SHAREDBUS_ADR_I[22] ), 
         .C(\SHAREDBUS_ADR_I[20] ), .D(\SHAREDBUS_ADR_I[16] ), .Z(n35796)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30634_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i30941_3_lut (.A(status_reg[0]), .B(inst1_FIFOfifo_rst), .C(n41345), 
         .Z(n36113)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30941_3_lut.init = 16'hcaca;
    LUT4 i30940_3_lut (.A(FIFOout_pins[0]), .B(inst3_Q[0]), .C(n41345), 
         .Z(n36112)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i30940_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_249 (.A(\SHAREDBUS_ADR_I[20] ), .B(n41347), 
         .C(n41303), .Z(n33894)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_3_lut_adj_249.init = 16'hfefe;
    LUT4 i1_2_lut_rep_885 (.A(\SHAREDBUS_ADR_I[27] ), .B(\SHAREDBUS_ADR_I[22] ), 
         .Z(n41290)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_885.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut_adj_250 (.A(\SHAREDBUS_ADR_I[27] ), .B(\SHAREDBUS_ADR_I[22] ), 
         .C(\SHAREDBUS_ADR_I[26] ), .D(\SHAREDBUS_ADR_I[29] ), .Z(n33784)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_250.init = 16'hfffe;
    LUT4 i1_4_lut_adj_251 (.A(n41246), .B(n33802), .C(n4865[18]), .D(n33720), 
         .Z(\FIFOwb_DAT_O[18] )) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_251.init = 16'hfffd;
    LUT4 i1_4_lut_adj_252 (.A(n41246), .B(n33802), .C(n4865[25]), .D(n33720), 
         .Z(\FIFOwb_DAT_O[25] )) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_252.init = 16'hfffd;
    PFUMX mux_1641_i32 (.BLUT(n1_adj_5866), .ALUT(n4865[31]), .C0(n37954), 
          .Z(\FIFOwb_DAT_O[31] ));
    PFUMX mux_1641_i31 (.BLUT(n1_adj_5865), .ALUT(n4865[30]), .C0(n37956), 
          .Z(\FIFOwb_DAT_O[30] ));
    PFUMX mux_1641_i28 (.BLUT(n1_adj_5864), .ALUT(n4865[27]), .C0(n37955), 
          .Z(\FIFOwb_DAT_O[27] ));
    PFUMX mux_1641_i27 (.BLUT(n1_adj_5863), .ALUT(n4865[26]), .C0(n37955), 
          .Z(\FIFOwb_DAT_O[26] ));
    PFUMX mux_1641_i24 (.BLUT(n1_adj_5862), .ALUT(n4865[23]), .C0(n37956), 
          .Z(\FIFOwb_DAT_O[23] ));
    PFUMX mux_1641_i21 (.BLUT(n1_adj_5861), .ALUT(n4865[20]), .C0(n37954), 
          .Z(\FIFOwb_DAT_O[20] ));
    PFUMX mux_1641_i20 (.BLUT(n1_adj_5860), .ALUT(n4865[19]), .C0(n37954), 
          .Z(\FIFOwb_DAT_O[19] ));
    PFUMX mux_1641_i17 (.BLUT(n1_adj_5859), .ALUT(n4865[16]), .C0(n37955), 
          .Z(\FIFOwb_DAT_O[16] ));
    PFUMX mux_1641_i11 (.BLUT(n1_adj_5858), .ALUT(n4865[10]), .C0(n37956), 
          .Z(\FIFOwb_DAT_O[10] ));
    PFUMX mux_1641_i9 (.BLUT(n1_adj_5857), .ALUT(n4865[8]), .C0(n37955), 
          .Z(\FIFOwb_DAT_O[8] ));
    PFUMX mux_1641_i6 (.BLUT(n1_adj_5856), .ALUT(n4865[5]), .C0(n37956), 
          .Z(\FIFOwb_DAT_O[5] ));
    PFUMX mux_1641_i2 (.BLUT(n36169), .ALUT(n36171), .C0(n37954), .Z(\FIFOwb_DAT_O[1] ));
    LUT4 i1_4_lut_adj_253 (.A(n41246), .B(n33802), .C(n4865[21]), .D(n33720), 
         .Z(\FIFOwb_DAT_O[21] )) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_253.init = 16'hfffd;
    LUT4 i1_4_lut_adj_254 (.A(n41246), .B(n33802), .C(n4865[28]), .D(n33720), 
         .Z(\FIFOwb_DAT_O[28] )) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_254.init = 16'hfffd;
    LUT4 i1_4_lut_adj_255 (.A(n41246), .B(n33802), .C(n4865[15]), .D(n33720), 
         .Z(\FIFOwb_DAT_O[15] )) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_255.init = 16'hfffd;
    LUT4 i1_4_lut_adj_256 (.A(n41246), .B(n33802), .C(n4865[13]), .D(n33720), 
         .Z(\FIFOwb_DAT_O[13] )) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_256.init = 16'hfffd;
    LUT4 i1_4_lut_adj_257 (.A(n41246), .B(n33802), .C(n4865[11]), .D(n33720), 
         .Z(\FIFOwb_DAT_O[11] )) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_257.init = 16'hfffd;
    LUT4 i1_4_lut_adj_258 (.A(n41246), .B(n33802), .C(n4865[9]), .D(n33720), 
         .Z(\FIFOwb_DAT_O[9] )) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_258.init = 16'hfffd;
    
endmodule
//
// Verilog Description of module fifo_dc_32x32
//

module fifo_dc_32x32 (inst3_Full, REF_CLK_c, inst1_FIFOfifo_rst, inst3_Empty, 
            GND_net, VCC_net, inst1_FIFOof_wr, inst1_FIFOif_rd, \SHAREDBUS_DAT_I[31] , 
            \SHAREDBUS_DAT_I[30] , \SHAREDBUS_DAT_I[29] , \SHAREDBUS_DAT_I[28] , 
            \SHAREDBUS_DAT_I[27] , \SHAREDBUS_DAT_I[26] , \SHAREDBUS_DAT_I[25] , 
            \SHAREDBUS_DAT_I[24] , n41343, n41342, n41341, n41340, 
            n41339, n41338, n41337, n41336, \SHAREDBUS_DAT_I[15] , 
            \SHAREDBUS_DAT_I[14] , \SHAREDBUS_DAT_I[13] , \SHAREDBUS_DAT_I[12] , 
            \SHAREDBUS_DAT_I[11] , \SHAREDBUS_DAT_I[10] , \SHAREDBUS_DAT_I[9] , 
            \SHAREDBUS_DAT_I[8] , n41335, n41334, n41333, n41332, 
            n41331, n41330, n41329, n41328, inst3_Q) /* synthesis NGD_DRC_MASK=1 */ ;
    output inst3_Full;
    input REF_CLK_c;
    input inst1_FIFOfifo_rst;
    output inst3_Empty;
    input GND_net;
    input VCC_net;
    input inst1_FIFOof_wr;
    input inst1_FIFOif_rd;
    input \SHAREDBUS_DAT_I[31] ;
    input \SHAREDBUS_DAT_I[30] ;
    input \SHAREDBUS_DAT_I[29] ;
    input \SHAREDBUS_DAT_I[28] ;
    input \SHAREDBUS_DAT_I[27] ;
    input \SHAREDBUS_DAT_I[26] ;
    input \SHAREDBUS_DAT_I[25] ;
    input \SHAREDBUS_DAT_I[24] ;
    input n41343;
    input n41342;
    input n41341;
    input n41340;
    input n41339;
    input n41338;
    input n41337;
    input n41336;
    input \SHAREDBUS_DAT_I[15] ;
    input \SHAREDBUS_DAT_I[14] ;
    input \SHAREDBUS_DAT_I[13] ;
    input \SHAREDBUS_DAT_I[12] ;
    input \SHAREDBUS_DAT_I[11] ;
    input \SHAREDBUS_DAT_I[10] ;
    input \SHAREDBUS_DAT_I[9] ;
    input \SHAREDBUS_DAT_I[8] ;
    input n41335;
    input n41334;
    input n41333;
    input n41332;
    input n41331;
    input n41330;
    input n41329;
    input n41328;
    output [31:0]inst3_Q;
    
    wire REF_CLK_c /* synthesis SET_AS_NETWORK=REF_CLK_c, is_clock=1 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(23[7:14])
    wire GND_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(23[7:15])
    wire VCC_net /* synthesis noprune=true */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/spi/fpgacfg.vhd(24[7:14])
    
    wire invout_1, iwcount_1, wren_i, wcount_1, iwcount_2, wcount_2, 
        iwcount_3, wcount_3, iwcount_4, wcount_4, iwcount_5, wcount_5, 
        w_gdata_0, w_gcount_0, w_gdata_1, w_gcount_1, w_gdata_2, w_gcount_2, 
        w_gdata_3, w_gcount_3, w_gdata_4, w_gcount_4, w_gcount_5, 
        wptr_0, wcount_0, wptr_1, wptr_2, wptr_3, wptr_4, wptr_5, 
        rRst, ircount_0, rden_i, rcount_0, ircount_1, rcount_1, 
        ircount_2, rcount_2, ircount_3, rcount_3, ircount_4, rcount_4, 
        ircount_5, rcount_5, r_gdata_0, r_gcount_0, r_gdata_1, r_gcount_1, 
        r_gdata_2, r_gcount_2, r_gdata_3, r_gcount_3, r_gdata_4, r_gcount_4, 
        r_gcount_5, rptr_0, rptr_1, rptr_2, rptr_3, rptr_4, rptr_5, 
        w_gcount_r0, w_gcount_r1, w_gcount_r2, w_gcount_r3, w_gcount_r4, 
        w_gcount_r5, r_gcount_w0, r_gcount_w1, r_gcount_w2, r_gcount_w3, 
        r_gcount_w4, r_gcount_w5, w_gcount_r20, w_gcount_r21, w_gcount_r22, 
        w_gcount_r23, w_gcount_r24, w_gcount_r25, r_gcount_w20, r_gcount_w21, 
        r_gcount_w22, r_gcount_w23, r_gcount_w24, r_gcount_w25, empty_d, 
        full_d, w_gctr_ci, iwcount_0, co0, co1, r_gctr_ci, co0_1, 
        co1_1, cmp_ci, wcount_r0, wcount_r1, co0_2, w_g2b_xor_cluster_0, 
        wcount_r3, co1_2, wcount_r4, empty_cmp_clr, empty_cmp_set, 
        empty_d_c, cmp_ci_1, rcount_w0, rcount_w1, co0_3, r_g2b_xor_cluster_0, 
        rcount_w3, co1_3, rcount_w4, full_cmp_clr, full_cmp_set, full_d_c, 
        invout_0;
    
    INV INV_1 (.A(inst3_Full), .Z(invout_1)) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    FD1P3DX FF_60 (.D(iwcount_1), .SP(wren_i), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(wcount_1)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(383[12:19])
    defparam FF_60.GSR = "ENABLED";
    FD1P3DX FF_59 (.D(iwcount_2), .SP(wren_i), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(wcount_2)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(387[12:19])
    defparam FF_59.GSR = "ENABLED";
    FD1P3DX FF_58 (.D(iwcount_3), .SP(wren_i), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(wcount_3)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(391[12:19])
    defparam FF_58.GSR = "ENABLED";
    FD1P3DX FF_57 (.D(iwcount_4), .SP(wren_i), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(wcount_4)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(395[12:19])
    defparam FF_57.GSR = "ENABLED";
    FD1P3DX FF_56 (.D(iwcount_5), .SP(wren_i), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(wcount_5)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(399[12:19])
    defparam FF_56.GSR = "ENABLED";
    FD1P3DX FF_55 (.D(w_gdata_0), .SP(wren_i), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_0)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(403[12:19])
    defparam FF_55.GSR = "ENABLED";
    FD1P3DX FF_54 (.D(w_gdata_1), .SP(wren_i), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_1)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(407[12:19])
    defparam FF_54.GSR = "ENABLED";
    FD1P3DX FF_53 (.D(w_gdata_2), .SP(wren_i), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_2)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(411[12:19])
    defparam FF_53.GSR = "ENABLED";
    FD1P3DX FF_52 (.D(w_gdata_3), .SP(wren_i), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_3)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(415[12:19])
    defparam FF_52.GSR = "ENABLED";
    FD1P3DX FF_51 (.D(w_gdata_4), .SP(wren_i), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_4)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(419[12:19])
    defparam FF_51.GSR = "ENABLED";
    FD1P3DX FF_50 (.D(wcount_5), .SP(wren_i), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_5)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(423[12:19])
    defparam FF_50.GSR = "ENABLED";
    FD1P3DX FF_49 (.D(wcount_0), .SP(wren_i), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(wptr_0)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(427[12:19])
    defparam FF_49.GSR = "ENABLED";
    FD1P3DX FF_48 (.D(wcount_1), .SP(wren_i), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(wptr_1)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(431[12:19])
    defparam FF_48.GSR = "ENABLED";
    FD1P3DX FF_47 (.D(wcount_2), .SP(wren_i), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(wptr_2)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(435[12:19])
    defparam FF_47.GSR = "ENABLED";
    FD1P3DX FF_46 (.D(wcount_3), .SP(wren_i), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(wptr_3)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(439[12:19])
    defparam FF_46.GSR = "ENABLED";
    FD1P3DX FF_45 (.D(wcount_4), .SP(wren_i), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(wptr_4)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(443[12:19])
    defparam FF_45.GSR = "ENABLED";
    FD1P3DX FF_44 (.D(wcount_5), .SP(wren_i), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(wptr_5)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(447[12:19])
    defparam FF_44.GSR = "ENABLED";
    FD1P3BX FF_43 (.D(ircount_0), .SP(rden_i), .CK(REF_CLK_c), .PD(rRst), 
            .Q(rcount_0)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(451[12:19])
    defparam FF_43.GSR = "ENABLED";
    FD1P3DX FF_42 (.D(ircount_1), .SP(rden_i), .CK(REF_CLK_c), .CD(rRst), 
            .Q(rcount_1)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(455[12:19])
    defparam FF_42.GSR = "ENABLED";
    FD1P3DX FF_41 (.D(ircount_2), .SP(rden_i), .CK(REF_CLK_c), .CD(rRst), 
            .Q(rcount_2)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(459[12:19])
    defparam FF_41.GSR = "ENABLED";
    FD1P3DX FF_40 (.D(ircount_3), .SP(rden_i), .CK(REF_CLK_c), .CD(rRst), 
            .Q(rcount_3)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(463[12:19])
    defparam FF_40.GSR = "ENABLED";
    FD1P3DX FF_39 (.D(ircount_4), .SP(rden_i), .CK(REF_CLK_c), .CD(rRst), 
            .Q(rcount_4)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(467[12:19])
    defparam FF_39.GSR = "ENABLED";
    FD1P3DX FF_38 (.D(ircount_5), .SP(rden_i), .CK(REF_CLK_c), .CD(rRst), 
            .Q(rcount_5)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(471[12:19])
    defparam FF_38.GSR = "ENABLED";
    FD1P3DX FF_37 (.D(r_gdata_0), .SP(rden_i), .CK(REF_CLK_c), .CD(rRst), 
            .Q(r_gcount_0)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(475[12:19])
    defparam FF_37.GSR = "ENABLED";
    FD1P3DX FF_36 (.D(r_gdata_1), .SP(rden_i), .CK(REF_CLK_c), .CD(rRst), 
            .Q(r_gcount_1)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(479[12:19])
    defparam FF_36.GSR = "ENABLED";
    FD1P3DX FF_35 (.D(r_gdata_2), .SP(rden_i), .CK(REF_CLK_c), .CD(rRst), 
            .Q(r_gcount_2)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(483[12:19])
    defparam FF_35.GSR = "ENABLED";
    FD1P3DX FF_34 (.D(r_gdata_3), .SP(rden_i), .CK(REF_CLK_c), .CD(rRst), 
            .Q(r_gcount_3)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(487[12:19])
    defparam FF_34.GSR = "ENABLED";
    FD1P3DX FF_33 (.D(r_gdata_4), .SP(rden_i), .CK(REF_CLK_c), .CD(rRst), 
            .Q(r_gcount_4)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(491[12:19])
    defparam FF_33.GSR = "ENABLED";
    FD1P3DX FF_32 (.D(rcount_5), .SP(rden_i), .CK(REF_CLK_c), .CD(rRst), 
            .Q(r_gcount_5)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(495[12:19])
    defparam FF_32.GSR = "ENABLED";
    FD1P3DX FF_31 (.D(rcount_0), .SP(rden_i), .CK(REF_CLK_c), .CD(rRst), 
            .Q(rptr_0)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(499[12:19])
    defparam FF_31.GSR = "ENABLED";
    FD1P3DX FF_30 (.D(rcount_1), .SP(rden_i), .CK(REF_CLK_c), .CD(rRst), 
            .Q(rptr_1)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(503[12:19])
    defparam FF_30.GSR = "ENABLED";
    FD1P3DX FF_29 (.D(rcount_2), .SP(rden_i), .CK(REF_CLK_c), .CD(rRst), 
            .Q(rptr_2)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(507[12:19])
    defparam FF_29.GSR = "ENABLED";
    FD1P3DX FF_28 (.D(rcount_3), .SP(rden_i), .CK(REF_CLK_c), .CD(rRst), 
            .Q(rptr_3)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(511[12:19])
    defparam FF_28.GSR = "ENABLED";
    FD1P3DX FF_27 (.D(rcount_4), .SP(rden_i), .CK(REF_CLK_c), .CD(rRst), 
            .Q(rptr_4)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(515[12:19])
    defparam FF_27.GSR = "ENABLED";
    FD1P3DX FF_26 (.D(rcount_5), .SP(rden_i), .CK(REF_CLK_c), .CD(rRst), 
            .Q(rptr_5)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(519[12:19])
    defparam FF_26.GSR = "ENABLED";
    FD1S3DX FF_25 (.D(w_gcount_0), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_r0)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(523[12:19])
    defparam FF_25.GSR = "ENABLED";
    FD1S3DX FF_24 (.D(w_gcount_1), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_r1)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(526[12:19])
    defparam FF_24.GSR = "ENABLED";
    FD1S3DX FF_23 (.D(w_gcount_2), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_r2)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(529[12:19])
    defparam FF_23.GSR = "ENABLED";
    FD1S3DX FF_22 (.D(w_gcount_3), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_r3)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(532[12:19])
    defparam FF_22.GSR = "ENABLED";
    FD1S3DX FF_21 (.D(w_gcount_4), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_r4)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(535[12:19])
    defparam FF_21.GSR = "ENABLED";
    FD1S3DX FF_20 (.D(w_gcount_5), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_r5)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(538[12:19])
    defparam FF_20.GSR = "ENABLED";
    FD1S3DX FF_19 (.D(r_gcount_0), .CK(REF_CLK_c), .CD(rRst), .Q(r_gcount_w0)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(541[12:19])
    defparam FF_19.GSR = "ENABLED";
    FD1S3DX FF_18 (.D(r_gcount_1), .CK(REF_CLK_c), .CD(rRst), .Q(r_gcount_w1)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(544[12:19])
    defparam FF_18.GSR = "ENABLED";
    FD1S3DX FF_17 (.D(r_gcount_2), .CK(REF_CLK_c), .CD(rRst), .Q(r_gcount_w2)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(547[12:19])
    defparam FF_17.GSR = "ENABLED";
    FD1S3DX FF_16 (.D(r_gcount_3), .CK(REF_CLK_c), .CD(rRst), .Q(r_gcount_w3)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(550[12:19])
    defparam FF_16.GSR = "ENABLED";
    FD1S3DX FF_15 (.D(r_gcount_4), .CK(REF_CLK_c), .CD(rRst), .Q(r_gcount_w4)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(553[12:19])
    defparam FF_15.GSR = "ENABLED";
    FD1S3DX FF_14 (.D(r_gcount_5), .CK(REF_CLK_c), .CD(rRst), .Q(r_gcount_w5)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(556[12:19])
    defparam FF_14.GSR = "ENABLED";
    FD1S3DX FF_13 (.D(w_gcount_r0), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_r20)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(559[12:19])
    defparam FF_13.GSR = "ENABLED";
    FD1S3DX FF_12 (.D(w_gcount_r1), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_r21)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(563[12:19])
    defparam FF_12.GSR = "ENABLED";
    FD1S3DX FF_11 (.D(w_gcount_r2), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_r22)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(567[12:19])
    defparam FF_11.GSR = "ENABLED";
    FD1S3DX FF_10 (.D(w_gcount_r3), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_r23)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(571[12:19])
    defparam FF_10.GSR = "ENABLED";
    FD1S3DX FF_9 (.D(w_gcount_r4), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_r24)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(575[11:18])
    defparam FF_9.GSR = "ENABLED";
    FD1S3DX FF_8 (.D(w_gcount_r5), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(w_gcount_r25)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(579[11:18])
    defparam FF_8.GSR = "ENABLED";
    FD1S3DX FF_7 (.D(r_gcount_w0), .CK(REF_CLK_c), .CD(rRst), .Q(r_gcount_w20)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(583[11:18])
    defparam FF_7.GSR = "ENABLED";
    FD1S3DX FF_6 (.D(r_gcount_w1), .CK(REF_CLK_c), .CD(rRst), .Q(r_gcount_w21)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(586[11:18])
    defparam FF_6.GSR = "ENABLED";
    FD1S3DX FF_5 (.D(r_gcount_w2), .CK(REF_CLK_c), .CD(rRst), .Q(r_gcount_w22)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(589[11:18])
    defparam FF_5.GSR = "ENABLED";
    FD1S3DX FF_4 (.D(r_gcount_w3), .CK(REF_CLK_c), .CD(rRst), .Q(r_gcount_w23)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(592[11:18])
    defparam FF_4.GSR = "ENABLED";
    FD1S3DX FF_3 (.D(r_gcount_w4), .CK(REF_CLK_c), .CD(rRst), .Q(r_gcount_w24)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(595[11:18])
    defparam FF_3.GSR = "ENABLED";
    FD1S3DX FF_2 (.D(r_gcount_w5), .CK(REF_CLK_c), .CD(rRst), .Q(r_gcount_w25)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(598[11:18])
    defparam FF_2.GSR = "ENABLED";
    FD1S3BX FF_1 (.D(empty_d), .CK(REF_CLK_c), .PD(rRst), .Q(inst3_Empty)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(601[11:18])
    defparam FF_1.GSR = "ENABLED";
    FD1S3DX FF_0 (.D(full_d), .CK(REF_CLK_c), .CD(inst1_FIFOfifo_rst), 
            .Q(inst3_Full)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(604[11:18])
    defparam FF_0.GSR = "ENABLED";
    CCU2C w_gctr_cia (.A0(GND_net), .B0(GND_net), .C0(VCC_net), .D0(VCC_net), 
          .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), .COUT(w_gctr_ci)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(607[17:22])
    defparam w_gctr_cia.INIT0 = 16'b0110011010101010;
    defparam w_gctr_cia.INIT1 = 16'b0110011010101010;
    defparam w_gctr_cia.INJECT1_0 = "NO";
    defparam w_gctr_cia.INJECT1_1 = "NO";
    CCU2C w_gctr_0 (.A0(wcount_0), .B0(GND_net), .C0(VCC_net), .D0(VCC_net), 
          .A1(wcount_1), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(w_gctr_ci), 
          .COUT(co0), .S0(iwcount_0), .S1(iwcount_1)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(614[15:20])
    defparam w_gctr_0.INIT0 = 16'b0110011010101010;
    defparam w_gctr_0.INIT1 = 16'b0110011010101010;
    defparam w_gctr_0.INJECT1_0 = "NO";
    defparam w_gctr_0.INJECT1_1 = "NO";
    CCU2C w_gctr_1 (.A0(wcount_2), .B0(GND_net), .C0(VCC_net), .D0(VCC_net), 
          .A1(wcount_3), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(co0), 
          .COUT(co1), .S0(iwcount_2), .S1(iwcount_3)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(622[15:20])
    defparam w_gctr_1.INIT0 = 16'b0110011010101010;
    defparam w_gctr_1.INIT1 = 16'b0110011010101010;
    defparam w_gctr_1.INJECT1_0 = "NO";
    defparam w_gctr_1.INJECT1_1 = "NO";
    CCU2C w_gctr_2 (.A0(wcount_4), .B0(GND_net), .C0(VCC_net), .D0(VCC_net), 
          .A1(wcount_5), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(co1), 
          .S0(iwcount_4), .S1(iwcount_5)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(630[15:20])
    defparam w_gctr_2.INIT0 = 16'b0110011010101010;
    defparam w_gctr_2.INIT1 = 16'b0110011010101010;
    defparam w_gctr_2.INJECT1_0 = "NO";
    defparam w_gctr_2.INJECT1_1 = "NO";
    CCU2C r_gctr_cia (.A0(GND_net), .B0(GND_net), .C0(VCC_net), .D0(VCC_net), 
          .A1(VCC_net), .B1(VCC_net), .C1(VCC_net), .D1(VCC_net), .COUT(r_gctr_ci)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(638[17:22])
    defparam r_gctr_cia.INIT0 = 16'b0110011010101010;
    defparam r_gctr_cia.INIT1 = 16'b0110011010101010;
    defparam r_gctr_cia.INJECT1_0 = "NO";
    defparam r_gctr_cia.INJECT1_1 = "NO";
    CCU2C r_gctr_0 (.A0(rcount_0), .B0(GND_net), .C0(VCC_net), .D0(VCC_net), 
          .A1(rcount_1), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(r_gctr_ci), 
          .COUT(co0_1), .S0(ircount_0), .S1(ircount_1)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(645[15:20])
    defparam r_gctr_0.INIT0 = 16'b0110011010101010;
    defparam r_gctr_0.INIT1 = 16'b0110011010101010;
    defparam r_gctr_0.INJECT1_0 = "NO";
    defparam r_gctr_0.INJECT1_1 = "NO";
    CCU2C r_gctr_1 (.A0(rcount_2), .B0(GND_net), .C0(VCC_net), .D0(VCC_net), 
          .A1(rcount_3), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(co0_1), 
          .COUT(co1_1), .S0(ircount_2), .S1(ircount_3)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(653[15:20])
    defparam r_gctr_1.INIT0 = 16'b0110011010101010;
    defparam r_gctr_1.INIT1 = 16'b0110011010101010;
    defparam r_gctr_1.INJECT1_0 = "NO";
    defparam r_gctr_1.INJECT1_1 = "NO";
    CCU2C r_gctr_2 (.A0(rcount_4), .B0(GND_net), .C0(VCC_net), .D0(VCC_net), 
          .A1(rcount_5), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(co1_1), 
          .S0(ircount_4), .S1(ircount_5)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(661[15:20])
    defparam r_gctr_2.INIT0 = 16'b0110011010101010;
    defparam r_gctr_2.INIT1 = 16'b0110011010101010;
    defparam r_gctr_2.INJECT1_0 = "NO";
    defparam r_gctr_2.INJECT1_1 = "NO";
    CCU2C empty_cmp_ci_a (.A0(GND_net), .B0(GND_net), .C0(VCC_net), .D0(VCC_net), 
          .A1(rden_i), .B1(rden_i), .C1(VCC_net), .D1(VCC_net), .COUT(cmp_ci)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(669[21:26])
    defparam empty_cmp_ci_a.INIT0 = 16'b0110011010101010;
    defparam empty_cmp_ci_a.INIT1 = 16'b0110011010101010;
    defparam empty_cmp_ci_a.INJECT1_0 = "NO";
    defparam empty_cmp_ci_a.INJECT1_1 = "NO";
    CCU2C empty_cmp_0 (.A0(rcount_0), .B0(wcount_r0), .C0(VCC_net), .D0(VCC_net), 
          .A1(rcount_1), .B1(wcount_r1), .C1(VCC_net), .D1(VCC_net), 
          .CIN(cmp_ci), .COUT(co0_2)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(676[18:23])
    defparam empty_cmp_0.INIT0 = 16'b1001100110101010;
    defparam empty_cmp_0.INIT1 = 16'b1001100110101010;
    defparam empty_cmp_0.INJECT1_0 = "NO";
    defparam empty_cmp_0.INJECT1_1 = "NO";
    CCU2C empty_cmp_1 (.A0(rcount_2), .B0(w_g2b_xor_cluster_0), .C0(VCC_net), 
          .D0(VCC_net), .A1(rcount_3), .B1(wcount_r3), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co0_2), .COUT(co1_2)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(683[18:23])
    defparam empty_cmp_1.INIT0 = 16'b1001100110101010;
    defparam empty_cmp_1.INIT1 = 16'b1001100110101010;
    defparam empty_cmp_1.INJECT1_0 = "NO";
    defparam empty_cmp_1.INJECT1_1 = "NO";
    CCU2C empty_cmp_2 (.A0(rcount_4), .B0(wcount_r4), .C0(VCC_net), .D0(VCC_net), 
          .A1(empty_cmp_set), .B1(empty_cmp_clr), .C1(VCC_net), .D1(VCC_net), 
          .CIN(co1_2), .COUT(empty_d_c)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(690[18:23])
    defparam empty_cmp_2.INIT0 = 16'b1001100110101010;
    defparam empty_cmp_2.INIT1 = 16'b1001100110101010;
    defparam empty_cmp_2.INJECT1_0 = "NO";
    defparam empty_cmp_2.INJECT1_1 = "NO";
    CCU2C a0 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(empty_d_c), 
          .S0(empty_d)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(698[9:14])
    defparam a0.INIT0 = 16'b0110011010101010;
    defparam a0.INIT1 = 16'b0110011010101010;
    defparam a0.INJECT1_0 = "NO";
    defparam a0.INJECT1_1 = "NO";
    CCU2C full_cmp_ci_a (.A0(GND_net), .B0(GND_net), .C0(VCC_net), .D0(VCC_net), 
          .A1(wren_i), .B1(wren_i), .C1(VCC_net), .D1(VCC_net), .COUT(cmp_ci_1)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(706[20:25])
    defparam full_cmp_ci_a.INIT0 = 16'b0110011010101010;
    defparam full_cmp_ci_a.INIT1 = 16'b0110011010101010;
    defparam full_cmp_ci_a.INJECT1_0 = "NO";
    defparam full_cmp_ci_a.INJECT1_1 = "NO";
    CCU2C full_cmp_0 (.A0(wcount_0), .B0(rcount_w0), .C0(VCC_net), .D0(VCC_net), 
          .A1(wcount_1), .B1(rcount_w1), .C1(VCC_net), .D1(VCC_net), 
          .CIN(cmp_ci_1), .COUT(co0_3)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(713[17:22])
    defparam full_cmp_0.INIT0 = 16'b1001100110101010;
    defparam full_cmp_0.INIT1 = 16'b1001100110101010;
    defparam full_cmp_0.INJECT1_0 = "NO";
    defparam full_cmp_0.INJECT1_1 = "NO";
    CCU2C full_cmp_1 (.A0(wcount_2), .B0(r_g2b_xor_cluster_0), .C0(VCC_net), 
          .D0(VCC_net), .A1(wcount_3), .B1(rcount_w3), .C1(VCC_net), 
          .D1(VCC_net), .CIN(co0_3), .COUT(co1_3)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(721[17:22])
    defparam full_cmp_1.INIT0 = 16'b1001100110101010;
    defparam full_cmp_1.INIT1 = 16'b1001100110101010;
    defparam full_cmp_1.INJECT1_0 = "NO";
    defparam full_cmp_1.INJECT1_1 = "NO";
    CCU2C full_cmp_2 (.A0(wcount_4), .B0(rcount_w4), .C0(VCC_net), .D0(VCC_net), 
          .A1(full_cmp_set), .B1(full_cmp_clr), .C1(VCC_net), .D1(VCC_net), 
          .CIN(co1_3), .COUT(full_d_c)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(728[17:22])
    defparam full_cmp_2.INIT0 = 16'b1001100110101010;
    defparam full_cmp_2.INIT1 = 16'b1001100110101010;
    defparam full_cmp_2.INJECT1_0 = "NO";
    defparam full_cmp_2.INJECT1_1 = "NO";
    CCU2C a1 (.A0(GND_net), .B0(GND_net), .C0(VCC_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(VCC_net), .D1(VCC_net), .CIN(full_d_c), 
          .S0(full_d)) /* synthesis syn_black_box=true, syn_unconnected_inputs="CIN", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(742[9:14])
    defparam a1.INIT0 = 16'b0110011010101010;
    defparam a1.INIT1 = 16'b0110011010101010;
    defparam a1.INJECT1_0 = "NO";
    defparam a1.INJECT1_1 = "NO";
    AND2 AND2_t12 (.A(inst1_FIFOof_wr), .B(invout_1), .Z(wren_i)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(226[15:19])
    AND2 AND2_t11 (.A(inst1_FIFOif_rd), .B(invout_0), .Z(rden_i)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(232[15:19])
    INV INV_0 (.A(inst3_Empty), .Z(invout_0)) /* synthesis LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    OR2 OR2_t10 (.A(inst1_FIFOfifo_rst), .B(inst1_FIFOfifo_rst), .Z(rRst)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(238[14:17])
    XOR2 XOR2_t9 (.A(wcount_0), .B(wcount_1), .Z(w_gdata_0)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(241[14:18])
    XOR2 XOR2_t8 (.A(wcount_1), .B(wcount_2), .Z(w_gdata_1)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(244[14:18])
    XOR2 XOR2_t7 (.A(wcount_2), .B(wcount_3), .Z(w_gdata_2)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(247[14:18])
    XOR2 XOR2_t6 (.A(wcount_3), .B(wcount_4), .Z(w_gdata_3)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(250[14:18])
    XOR2 XOR2_t5 (.A(wcount_4), .B(wcount_5), .Z(w_gdata_4)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(253[14:18])
    XOR2 XOR2_t4 (.A(rcount_0), .B(rcount_1), .Z(r_gdata_0)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(256[14:18])
    XOR2 XOR2_t3 (.A(rcount_1), .B(rcount_2), .Z(r_gdata_1)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(259[14:18])
    XOR2 XOR2_t2 (.A(rcount_2), .B(rcount_3), .Z(r_gdata_2)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(262[14:18])
    XOR2 XOR2_t1 (.A(rcount_3), .B(rcount_4), .Z(r_gdata_3)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(265[14:18])
    XOR2 XOR2_t0 (.A(rcount_4), .B(rcount_5), .Z(r_gdata_4)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(268[14:18])
    ROM16X1A LUT4_13 (.AD0(w_gcount_r25), .AD1(w_gcount_r24), .AD2(w_gcount_r23), 
            .AD3(w_gcount_r22), .DO0(w_g2b_xor_cluster_0)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    defparam LUT4_13.initval = 16'b0110100110010110;
    ROM16X1A LUT4_12 (.AD0(GND_net), .AD1(GND_net), .AD2(w_gcount_r25), 
            .AD3(w_gcount_r24), .DO0(wcount_r4)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    defparam LUT4_12.initval = 16'b0110100110010110;
    ROM16X1A LUT4_11 (.AD0(GND_net), .AD1(w_gcount_r25), .AD2(w_gcount_r24), 
            .AD3(w_gcount_r23), .DO0(wcount_r3)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    defparam LUT4_11.initval = 16'b0110100110010110;
    ROM16X1A LUT4_10 (.AD0(wcount_r4), .AD1(w_gcount_r23), .AD2(w_gcount_r22), 
            .AD3(w_gcount_r21), .DO0(wcount_r1)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    defparam LUT4_10.initval = 16'b0110100110010110;
    ROM16X1A LUT4_9 (.AD0(wcount_r3), .AD1(w_gcount_r22), .AD2(w_gcount_r21), 
            .AD3(w_gcount_r20), .DO0(wcount_r0)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    defparam LUT4_9.initval = 16'b0110100110010110;
    ROM16X1A LUT4_8 (.AD0(r_gcount_w25), .AD1(r_gcount_w24), .AD2(r_gcount_w23), 
            .AD3(r_gcount_w22), .DO0(r_g2b_xor_cluster_0)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    defparam LUT4_8.initval = 16'b0110100110010110;
    ROM16X1A LUT4_7 (.AD0(GND_net), .AD1(GND_net), .AD2(r_gcount_w25), 
            .AD3(r_gcount_w24), .DO0(rcount_w4)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    defparam LUT4_7.initval = 16'b0110100110010110;
    ROM16X1A LUT4_6 (.AD0(GND_net), .AD1(r_gcount_w25), .AD2(r_gcount_w24), 
            .AD3(r_gcount_w23), .DO0(rcount_w3)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    defparam LUT4_6.initval = 16'b0110100110010110;
    ROM16X1A LUT4_5 (.AD0(rcount_w4), .AD1(r_gcount_w23), .AD2(r_gcount_w22), 
            .AD3(r_gcount_w21), .DO0(rcount_w1)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    defparam LUT4_5.initval = 16'b0110100110010110;
    ROM16X1A LUT4_4 (.AD0(rcount_w3), .AD1(r_gcount_w22), .AD2(r_gcount_w21), 
            .AD3(r_gcount_w20), .DO0(rcount_w0)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    defparam LUT4_4.initval = 16'b0110100110010110;
    ROM16X1A LUT4_3 (.AD0(GND_net), .AD1(w_gcount_r25), .AD2(rcount_5), 
            .AD3(rptr_5), .DO0(empty_cmp_set)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    defparam LUT4_3.initval = 16'b0000010000010000;
    ROM16X1A LUT4_2 (.AD0(GND_net), .AD1(w_gcount_r25), .AD2(rcount_5), 
            .AD3(rptr_5), .DO0(empty_cmp_clr)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    defparam LUT4_2.initval = 16'b0001000000000100;
    ROM16X1A LUT4_1 (.AD0(GND_net), .AD1(r_gcount_w25), .AD2(wcount_5), 
            .AD3(wptr_5), .DO0(full_cmp_set)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    defparam LUT4_1.initval = 16'b0000000101000000;
    ROM16X1A LUT4_0 (.AD0(GND_net), .AD1(r_gcount_w25), .AD2(wcount_5), 
            .AD3(wptr_5), .DO0(full_cmp_clr)) /* synthesis syn_black_box=true, syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    defparam LUT4_0.initval = 16'b0100000000000001;
    PDPW16KD pdp_ram_0_0_0 (.DI0(n41328), .DI1(n41329), .DI2(n41330), 
            .DI3(n41331), .DI4(n41332), .DI5(n41333), .DI6(n41334), 
            .DI7(n41335), .DI8(\SHAREDBUS_DAT_I[8] ), .DI9(\SHAREDBUS_DAT_I[9] ), 
            .DI10(\SHAREDBUS_DAT_I[10] ), .DI11(\SHAREDBUS_DAT_I[11] ), 
            .DI12(\SHAREDBUS_DAT_I[12] ), .DI13(\SHAREDBUS_DAT_I[13] ), 
            .DI14(\SHAREDBUS_DAT_I[14] ), .DI15(\SHAREDBUS_DAT_I[15] ), 
            .DI16(n41336), .DI17(n41337), .DI18(n41338), .DI19(n41339), 
            .DI20(n41340), .DI21(n41341), .DI22(n41342), .DI23(n41343), 
            .DI24(\SHAREDBUS_DAT_I[24] ), .DI25(\SHAREDBUS_DAT_I[25] ), 
            .DI26(\SHAREDBUS_DAT_I[26] ), .DI27(\SHAREDBUS_DAT_I[27] ), 
            .DI28(\SHAREDBUS_DAT_I[28] ), .DI29(\SHAREDBUS_DAT_I[29] ), 
            .DI30(\SHAREDBUS_DAT_I[30] ), .DI31(\SHAREDBUS_DAT_I[31] ), 
            .DI32(GND_net), .DI33(GND_net), .DI34(GND_net), .DI35(GND_net), 
            .ADW0(wptr_0), .ADW1(wptr_1), .ADW2(wptr_2), .ADW3(wptr_3), 
            .ADW4(wptr_4), .ADW5(GND_net), .ADW6(GND_net), .ADW7(GND_net), 
            .ADW8(GND_net), .BE0(VCC_net), .BE1(VCC_net), .BE2(VCC_net), 
            .BE3(VCC_net), .CEW(wren_i), .CLKW(REF_CLK_c), .CSW0(VCC_net), 
            .CSW1(GND_net), .CSW2(GND_net), .ADR0(GND_net), .ADR1(GND_net), 
            .ADR2(GND_net), .ADR3(GND_net), .ADR4(GND_net), .ADR5(rptr_0), 
            .ADR6(rptr_1), .ADR7(rptr_2), .ADR8(rptr_3), .ADR9(rptr_4), 
            .ADR10(GND_net), .ADR11(GND_net), .ADR12(GND_net), .ADR13(GND_net), 
            .CER(rden_i), .OCER(rden_i), .CLKR(REF_CLK_c), .CSR0(GND_net), 
            .CSR1(GND_net), .CSR2(GND_net), .RST(inst1_FIFOfifo_rst), 
            .DO0(inst3_Q[18]), .DO1(inst3_Q[19]), .DO2(inst3_Q[20]), .DO3(inst3_Q[21]), 
            .DO4(inst3_Q[22]), .DO5(inst3_Q[23]), .DO6(inst3_Q[24]), .DO7(inst3_Q[25]), 
            .DO8(inst3_Q[26]), .DO9(inst3_Q[27]), .DO10(inst3_Q[28]), 
            .DO11(inst3_Q[29]), .DO12(inst3_Q[30]), .DO13(inst3_Q[31]), 
            .DO18(inst3_Q[0]), .DO19(inst3_Q[1]), .DO20(inst3_Q[2]), .DO21(inst3_Q[3]), 
            .DO22(inst3_Q[4]), .DO23(inst3_Q[5]), .DO24(inst3_Q[6]), .DO25(inst3_Q[7]), 
            .DO26(inst3_Q[8]), .DO27(inst3_Q[9]), .DO28(inst3_Q[10]), 
            .DO29(inst3_Q[11]), .DO30(inst3_Q[12]), .DO31(inst3_Q[13]), 
            .DO32(inst3_Q[14]), .DO33(inst3_Q[15]), .DO34(inst3_Q[16]), 
            .DO35(inst3_Q[17])) /* synthesis syn_black_box=true, MEM_LPC_FILE="fifo_dc_32x32.lpc", MEM_INIT_FILE="", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/src/top.vhd(138[9:34])
    defparam pdp_ram_0_0_0.DATA_WIDTH_W = 36;
    defparam pdp_ram_0_0_0.DATA_WIDTH_R = 36;
    defparam pdp_ram_0_0_0.GSR = "ENABLED";
    defparam pdp_ram_0_0_0.REGMODE = "NOREG";
    defparam pdp_ram_0_0_0.RESETMODE = "ASYNC";
    defparam pdp_ram_0_0_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam pdp_ram_0_0_0.CSDECODE_W = "0b001";
    defparam pdp_ram_0_0_0.CSDECODE_R = "0b000";
    defparam pdp_ram_0_0_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam pdp_ram_0_0_0.INIT_DATA = "STATIC";
    FD1P3BX FF_61 (.D(iwcount_0), .SP(wren_i), .CK(REF_CLK_c), .PD(inst1_FIFOfifo_rst), 
            .Q(wcount_0)) /* synthesis syn_black_box=true, GSR="ENABLED", syn_instantiated=1, LSE_LINE_FILE_ID=61, LSE_LCOL=9, LSE_RCOL=34, LSE_LLINE=138, LSE_RLINE=138 */ ;   // d:/darbas/lattice/orange_crab/lm32_tutor/ip/fifo_dc_32x32/fifo_dc_32x32/fifo_dc_32x32.vhd(379[12:19])
    defparam FF_61.GSR = "ENABLED";
    
endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.12.1.454 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.12/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch sa5p00 -type bram -wp 10 -rp 0011 -data_width 32 -num_rows 8192 -rdata_width 32 -gsr ENABLED -sync_reset -memformat hex -cascade -1 -n pmi_ram_dpEhnonessen321381923213819211e08d7f -pmi -lang verilog  */
/* Sun Jan 23 21:09:14 2022 */


`timescale 1 ns / 1 ps
module pmi_ram_dpEhnonessen321381923213819211e08d7f (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [12:0] WrAddress;
    input wire [12:0] RdAddress;
    input wire [31:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [31:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[1]), 
        .DIA0(Data[0]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[1]), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[3]), 
        .DIA0(Data[2]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[3]), .DOB0(Q[2]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[5]), 
        .DIA0(Data[4]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[5]), .DOB0(Q[4]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[7]), 
        .DIA0(Data[6]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[7]), .DOB0(Q[6]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[9]), 
        .DIA0(Data[8]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[9]), .DOB0(Q[8]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[11]), 
        .DIA0(Data[10]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[11]), .DOB0(Q[10]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[13]), 
        .DIA0(Data[12]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[13]), .DOB0(Q[12]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[15]), 
        .DIA0(Data[14]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[15]), .DOB0(Q[14]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[17]), 
        .DIA0(Data[16]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[17]), .DOB0(Q[16]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[19]), 
        .DIA0(Data[18]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[19]), .DOB0(Q[18]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[21]), 
        .DIA0(Data[20]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[21]), .DOB0(Q[20]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[23]), 
        .DIA0(Data[22]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[23]), .DOB0(Q[22]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[25]), 
        .DIA0(Data[24]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[25]), .DOB0(Q[24]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[27]), 
        .DIA0(Data[26]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[27]), .DOB0(Q[26]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[29]), 
        .DIA0(Data[28]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[29]), .DOB0(Q[28]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[31]), 
        .DIA0(Data[30]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[31]), .DOB0(Q[30]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.12.1.454 */
/* Module Version: 3.5 */
/* C:/lscc/diamond/3.12/ispfpga/bin/nt64/scuba -w -arch sa5p00 -n pmi_addsubEo3232491b9e8 -bb -bus_exp 7 -type addsub -width 32 -unsigned -port ci -port co -pmi -lang verilog  */
/* Sun Jan 23 21:09:14 2022 */


`timescale 1 ns / 1 ps
module pmi_addsubEo3232491b9e8 (DataA, DataB, Cin, Add_Sub, Result, Cout, 
    Overflow)/* synthesis NGD_DRC_MASK=1 */;
    input wire [31:0] DataA;
    input wire [31:0] DataB;
    input wire Cin;
    input wire Add_Sub;
    output wire [31:0] Result;
    output wire Cout;
    output wire Overflow;

    wire ci_k;
    wire precin;
    wire co0;
    wire co1;
    wire co2;
    wire co3;
    wire co4;
    wire co5;
    wire co6;
    wire co7;
    wire co8;
    wire co9;
    wire co10;
    wire co11;
    wire co12;
    wire co13;
    wire co14;
    wire add_sub_inv;
    wire co15;
    wire co16d;
    wire scuba_vhi;
    wire scuba_vlo;
    wire co16;

    XNOR2 XNOR2_t0 (.A(Cin), .B(Add_Sub), .Z(ci_k));

    INV INV_0 (.A(Add_Sub), .Z(add_sub_inv));

    defparam precin_inst102.INJECT1_1 = "NO" ;
    defparam precin_inst102.INJECT1_0 = "NO" ;
    defparam precin_inst102.INIT1 =  16'h0000 ;
    defparam precin_inst102.INIT0 =  16'h0000 ;
    CCU2C precin_inst102 (.A0(scuba_vhi), .A1(scuba_vhi), .B0(scuba_vhi), 
        .B1(scuba_vhi), .C0(scuba_vhi), .C1(scuba_vhi), .D0(scuba_vhi), 
        .D1(scuba_vhi), .CIN(), .S0(), .S1(), .COUT(precin));

    defparam addsub_0.INJECT1_1 = "NO" ;
    defparam addsub_0.INJECT1_0 = "NO" ;
    defparam addsub_0.INIT1 =  16'h69AA ;
    defparam addsub_0.INIT0 =  16'h69AA ;
    CCU2C addsub_0 (.A0(Cin), .A1(DataA[0]), .B0(ci_k), .B1(DataB[0]), .C0(Add_Sub), 
        .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(precin), .S0(), 
        .S1(Result[0]), .COUT(co0));

    defparam addsub_1.INJECT1_1 = "NO" ;
    defparam addsub_1.INJECT1_0 = "NO" ;
    defparam addsub_1.INIT1 =  16'h69AA ;
    defparam addsub_1.INIT0 =  16'h69AA ;
    CCU2C addsub_1 (.A0(DataA[1]), .A1(DataA[2]), .B0(DataB[1]), .B1(DataB[2]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co0), 
        .S0(Result[1]), .S1(Result[2]), .COUT(co1));

    defparam addsub_2.INJECT1_1 = "NO" ;
    defparam addsub_2.INJECT1_0 = "NO" ;
    defparam addsub_2.INIT1 =  16'h69AA ;
    defparam addsub_2.INIT0 =  16'h69AA ;
    CCU2C addsub_2 (.A0(DataA[3]), .A1(DataA[4]), .B0(DataB[3]), .B1(DataB[4]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co1), 
        .S0(Result[3]), .S1(Result[4]), .COUT(co2));

    defparam addsub_3.INJECT1_1 = "NO" ;
    defparam addsub_3.INJECT1_0 = "NO" ;
    defparam addsub_3.INIT1 =  16'h69AA ;
    defparam addsub_3.INIT0 =  16'h69AA ;
    CCU2C addsub_3 (.A0(DataA[5]), .A1(DataA[6]), .B0(DataB[5]), .B1(DataB[6]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co2), 
        .S0(Result[5]), .S1(Result[6]), .COUT(co3));

    defparam addsub_4.INJECT1_1 = "NO" ;
    defparam addsub_4.INJECT1_0 = "NO" ;
    defparam addsub_4.INIT1 =  16'h69AA ;
    defparam addsub_4.INIT0 =  16'h69AA ;
    CCU2C addsub_4 (.A0(DataA[7]), .A1(DataA[8]), .B0(DataB[7]), .B1(DataB[8]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co3), 
        .S0(Result[7]), .S1(Result[8]), .COUT(co4));

    defparam addsub_5.INJECT1_1 = "NO" ;
    defparam addsub_5.INJECT1_0 = "NO" ;
    defparam addsub_5.INIT1 =  16'h69AA ;
    defparam addsub_5.INIT0 =  16'h69AA ;
    CCU2C addsub_5 (.A0(DataA[9]), .A1(DataA[10]), .B0(DataB[9]), .B1(DataB[10]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co4), 
        .S0(Result[9]), .S1(Result[10]), .COUT(co5));

    defparam addsub_6.INJECT1_1 = "NO" ;
    defparam addsub_6.INJECT1_0 = "NO" ;
    defparam addsub_6.INIT1 =  16'h69AA ;
    defparam addsub_6.INIT0 =  16'h69AA ;
    CCU2C addsub_6 (.A0(DataA[11]), .A1(DataA[12]), .B0(DataB[11]), .B1(DataB[12]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co5), 
        .S0(Result[11]), .S1(Result[12]), .COUT(co6));

    defparam addsub_7.INJECT1_1 = "NO" ;
    defparam addsub_7.INJECT1_0 = "NO" ;
    defparam addsub_7.INIT1 =  16'h69AA ;
    defparam addsub_7.INIT0 =  16'h69AA ;
    CCU2C addsub_7 (.A0(DataA[13]), .A1(DataA[14]), .B0(DataB[13]), .B1(DataB[14]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co6), 
        .S0(Result[13]), .S1(Result[14]), .COUT(co7));

    defparam addsub_8.INJECT1_1 = "NO" ;
    defparam addsub_8.INJECT1_0 = "NO" ;
    defparam addsub_8.INIT1 =  16'h69AA ;
    defparam addsub_8.INIT0 =  16'h69AA ;
    CCU2C addsub_8 (.A0(DataA[15]), .A1(DataA[16]), .B0(DataB[15]), .B1(DataB[16]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co7), 
        .S0(Result[15]), .S1(Result[16]), .COUT(co8));

    defparam addsub_9.INJECT1_1 = "NO" ;
    defparam addsub_9.INJECT1_0 = "NO" ;
    defparam addsub_9.INIT1 =  16'h69AA ;
    defparam addsub_9.INIT0 =  16'h69AA ;
    CCU2C addsub_9 (.A0(DataA[17]), .A1(DataA[18]), .B0(DataB[17]), .B1(DataB[18]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co8), 
        .S0(Result[17]), .S1(Result[18]), .COUT(co9));

    defparam addsub_10.INJECT1_1 = "NO" ;
    defparam addsub_10.INJECT1_0 = "NO" ;
    defparam addsub_10.INIT1 =  16'h69AA ;
    defparam addsub_10.INIT0 =  16'h69AA ;
    CCU2C addsub_10 (.A0(DataA[19]), .A1(DataA[20]), .B0(DataB[19]), .B1(DataB[20]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co9), 
        .S0(Result[19]), .S1(Result[20]), .COUT(co10));

    defparam addsub_11.INJECT1_1 = "NO" ;
    defparam addsub_11.INJECT1_0 = "NO" ;
    defparam addsub_11.INIT1 =  16'h69AA ;
    defparam addsub_11.INIT0 =  16'h69AA ;
    CCU2C addsub_11 (.A0(DataA[21]), .A1(DataA[22]), .B0(DataB[21]), .B1(DataB[22]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co10), 
        .S0(Result[21]), .S1(Result[22]), .COUT(co11));

    defparam addsub_12.INJECT1_1 = "NO" ;
    defparam addsub_12.INJECT1_0 = "NO" ;
    defparam addsub_12.INIT1 =  16'h69AA ;
    defparam addsub_12.INIT0 =  16'h69AA ;
    CCU2C addsub_12 (.A0(DataA[23]), .A1(DataA[24]), .B0(DataB[23]), .B1(DataB[24]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co11), 
        .S0(Result[23]), .S1(Result[24]), .COUT(co12));

    defparam addsub_13.INJECT1_1 = "NO" ;
    defparam addsub_13.INJECT1_0 = "NO" ;
    defparam addsub_13.INIT1 =  16'h69AA ;
    defparam addsub_13.INIT0 =  16'h69AA ;
    CCU2C addsub_13 (.A0(DataA[25]), .A1(DataA[26]), .B0(DataB[25]), .B1(DataB[26]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co12), 
        .S0(Result[25]), .S1(Result[26]), .COUT(co13));

    defparam addsub_14.INJECT1_1 = "NO" ;
    defparam addsub_14.INJECT1_0 = "NO" ;
    defparam addsub_14.INIT1 =  16'h69AA ;
    defparam addsub_14.INIT0 =  16'h69AA ;
    CCU2C addsub_14 (.A0(DataA[27]), .A1(DataA[28]), .B0(DataB[27]), .B1(DataB[28]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co13), 
        .S0(Result[27]), .S1(Result[28]), .COUT(co14));

    defparam addsub_15.INJECT1_1 = "NO" ;
    defparam addsub_15.INJECT1_0 = "NO" ;
    defparam addsub_15.INIT1 =  16'h69AA ;
    defparam addsub_15.INIT0 =  16'h69AA ;
    CCU2C addsub_15 (.A0(DataA[29]), .A1(DataA[30]), .B0(DataB[29]), .B1(DataB[30]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co14), 
        .S0(Result[29]), .S1(Result[30]), .COUT(co15));

    defparam addsub_16.INJECT1_1 = "NO" ;
    defparam addsub_16.INJECT1_0 = "NO" ;
    defparam addsub_16.INIT1 =  16'h69AA ;
    defparam addsub_16.INIT0 =  16'h69AA ;
    CCU2C addsub_16 (.A0(DataA[31]), .A1(scuba_vlo), .B0(DataB[31]), .B1(add_sub_inv), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co15), 
        .S0(Result[31]), .S1(Cout), .COUT(co16));

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam addsubd.INJECT1_1 = "NO" ;
    defparam addsubd.INJECT1_0 = "NO" ;
    defparam addsubd.INIT1 =  16'h66AA ;
    defparam addsubd.INIT0 =  16'h66AA ;
    CCU2C addsubd (.A0(scuba_vlo), .A1(scuba_vlo), .B0(scuba_vlo), .B1(scuba_vlo), 
        .C0(scuba_vhi), .C1(scuba_vhi), .D0(scuba_vhi), .D1(scuba_vhi), 
        .CIN(co16), .S0(co16d), .S1(), .COUT());



    // exemplar begin
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.12.1.454 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.12/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch sa5p00 -type bram -wp 10 -rp 0011 -data_width 32 -num_rows 8192 -rdata_width 32 -gsr ENABLED -sync_reset -memformat hex -cascade -1 -n pmi_ram_dpEhnonessen321381923213819211e08d7f -pmi -lang verilog  */
/* Sun Feb 06 15:10:23 2022 */


`timescale 1 ns / 1 ps
module pmi_ram_dpEhnonessen321381923213819211e08d7f (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [12:0] WrAddress;
    input wire [12:0] RdAddress;
    input wire [31:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [31:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[1]), 
        .DIA0(Data[0]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[1]), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[3]), 
        .DIA0(Data[2]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[3]), .DOB0(Q[2]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[5]), 
        .DIA0(Data[4]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[5]), .DOB0(Q[4]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[7]), 
        .DIA0(Data[6]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[7]), .DOB0(Q[6]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[9]), 
        .DIA0(Data[8]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[9]), .DOB0(Q[8]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[11]), 
        .DIA0(Data[10]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[11]), .DOB0(Q[10]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[13]), 
        .DIA0(Data[12]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[13]), .DOB0(Q[12]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[15]), 
        .DIA0(Data[14]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[15]), .DOB0(Q[14]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[17]), 
        .DIA0(Data[16]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[17]), .DOB0(Q[16]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[19]), 
        .DIA0(Data[18]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[19]), .DOB0(Q[18]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[21]), 
        .DIA0(Data[20]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[21]), .DOB0(Q[20]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[23]), 
        .DIA0(Data[22]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[23]), .DOB0(Q[22]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[25]), 
        .DIA0(Data[24]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[25]), .DOB0(Q[24]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[27]), 
        .DIA0(Data[26]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[27]), .DOB0(Q[26]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[29]), 
        .DIA0(Data[28]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[29]), .DOB0(Q[28]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.RESETMODE = "SYNC" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.REGMODE_B = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.REGMODE_A = "NOREG" ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.DATA_WIDTH_B = 2 ;
    defparam pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0.DATA_WIDTH_A = 2 ;
    DP16KD pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(Data[31]), 
        .DIA0(Data[30]), .ADA13(WrAddress[12]), .ADA12(WrAddress[11]), .ADA11(WrAddress[10]), 
        .ADA10(WrAddress[9]), .ADA9(WrAddress[8]), .ADA8(WrAddress[7]), 
        .ADA7(WrAddress[6]), .ADA6(WrAddress[5]), .ADA5(WrAddress[4]), .ADA4(WrAddress[3]), 
        .ADA3(WrAddress[2]), .ADA2(WrAddress[1]), .ADA1(WrAddress[0]), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[12]), .ADB12(RdAddress[11]), 
        .ADB11(RdAddress[10]), .ADB10(RdAddress[9]), .ADB9(RdAddress[8]), 
        .ADB8(RdAddress[7]), .ADB7(RdAddress[6]), .ADB6(RdAddress[5]), .ADB5(RdAddress[4]), 
        .ADB4(RdAddress[3]), .ADB3(RdAddress[2]), .ADB2(RdAddress[1]), .ADB1(RdAddress[0]), 
        .ADB0(scuba_vlo), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), 
        .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), 
        .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(Q[31]), .DOB0(Q[30]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_0_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_1_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_2_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_3_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_4_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_5_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_6_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_7_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_8_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_9_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_10_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_11_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_12_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_13_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_14_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0 MEM_LPC_FILE pmi_ram_dpEhnonessen321381923213819211e08d7f__PMIP__8192__32__32H
    // exemplar attribute pmi_ram_dpEhnonessen321381923213819211e08d7f_0_15_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.12.1.454 */
/* Module Version: 3.5 */
/* C:/lscc/diamond/3.12/ispfpga/bin/nt64/scuba -w -arch sa5p00 -n pmi_addsubEo3232491b9e8 -bb -bus_exp 7 -type addsub -width 32 -unsigned -port ci -port co -pmi -lang verilog  */
/* Sun Feb 06 15:10:23 2022 */


`timescale 1 ns / 1 ps
module pmi_addsubEo3232491b9e8 (DataA, DataB, Cin, Add_Sub, Result, Cout, 
    Overflow)/* synthesis NGD_DRC_MASK=1 */;
    input wire [31:0] DataA;
    input wire [31:0] DataB;
    input wire Cin;
    input wire Add_Sub;
    output wire [31:0] Result;
    output wire Cout;
    output wire Overflow;

    wire ci_k;
    wire precin;
    wire co0;
    wire co1;
    wire co2;
    wire co3;
    wire co4;
    wire co5;
    wire co6;
    wire co7;
    wire co8;
    wire co9;
    wire co10;
    wire co11;
    wire co12;
    wire co13;
    wire co14;
    wire add_sub_inv;
    wire co15;
    wire co16d;
    wire scuba_vhi;
    wire scuba_vlo;
    wire co16;

    XNOR2 XNOR2_t0 (.A(Cin), .B(Add_Sub), .Z(ci_k));

    INV INV_0 (.A(Add_Sub), .Z(add_sub_inv));

    defparam precin_inst102.INJECT1_1 = "NO" ;
    defparam precin_inst102.INJECT1_0 = "NO" ;
    defparam precin_inst102.INIT1 =  16'h0000 ;
    defparam precin_inst102.INIT0 =  16'h0000 ;
    CCU2C precin_inst102 (.A0(scuba_vhi), .A1(scuba_vhi), .B0(scuba_vhi), 
        .B1(scuba_vhi), .C0(scuba_vhi), .C1(scuba_vhi), .D0(scuba_vhi), 
        .D1(scuba_vhi), .CIN(), .S0(), .S1(), .COUT(precin));

    defparam addsub_0.INJECT1_1 = "NO" ;
    defparam addsub_0.INJECT1_0 = "NO" ;
    defparam addsub_0.INIT1 =  16'h69AA ;
    defparam addsub_0.INIT0 =  16'h69AA ;
    CCU2C addsub_0 (.A0(Cin), .A1(DataA[0]), .B0(ci_k), .B1(DataB[0]), .C0(Add_Sub), 
        .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(precin), .S0(), 
        .S1(Result[0]), .COUT(co0));

    defparam addsub_1.INJECT1_1 = "NO" ;
    defparam addsub_1.INJECT1_0 = "NO" ;
    defparam addsub_1.INIT1 =  16'h69AA ;
    defparam addsub_1.INIT0 =  16'h69AA ;
    CCU2C addsub_1 (.A0(DataA[1]), .A1(DataA[2]), .B0(DataB[1]), .B1(DataB[2]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co0), 
        .S0(Result[1]), .S1(Result[2]), .COUT(co1));

    defparam addsub_2.INJECT1_1 = "NO" ;
    defparam addsub_2.INJECT1_0 = "NO" ;
    defparam addsub_2.INIT1 =  16'h69AA ;
    defparam addsub_2.INIT0 =  16'h69AA ;
    CCU2C addsub_2 (.A0(DataA[3]), .A1(DataA[4]), .B0(DataB[3]), .B1(DataB[4]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co1), 
        .S0(Result[3]), .S1(Result[4]), .COUT(co2));

    defparam addsub_3.INJECT1_1 = "NO" ;
    defparam addsub_3.INJECT1_0 = "NO" ;
    defparam addsub_3.INIT1 =  16'h69AA ;
    defparam addsub_3.INIT0 =  16'h69AA ;
    CCU2C addsub_3 (.A0(DataA[5]), .A1(DataA[6]), .B0(DataB[5]), .B1(DataB[6]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co2), 
        .S0(Result[5]), .S1(Result[6]), .COUT(co3));

    defparam addsub_4.INJECT1_1 = "NO" ;
    defparam addsub_4.INJECT1_0 = "NO" ;
    defparam addsub_4.INIT1 =  16'h69AA ;
    defparam addsub_4.INIT0 =  16'h69AA ;
    CCU2C addsub_4 (.A0(DataA[7]), .A1(DataA[8]), .B0(DataB[7]), .B1(DataB[8]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co3), 
        .S0(Result[7]), .S1(Result[8]), .COUT(co4));

    defparam addsub_5.INJECT1_1 = "NO" ;
    defparam addsub_5.INJECT1_0 = "NO" ;
    defparam addsub_5.INIT1 =  16'h69AA ;
    defparam addsub_5.INIT0 =  16'h69AA ;
    CCU2C addsub_5 (.A0(DataA[9]), .A1(DataA[10]), .B0(DataB[9]), .B1(DataB[10]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co4), 
        .S0(Result[9]), .S1(Result[10]), .COUT(co5));

    defparam addsub_6.INJECT1_1 = "NO" ;
    defparam addsub_6.INJECT1_0 = "NO" ;
    defparam addsub_6.INIT1 =  16'h69AA ;
    defparam addsub_6.INIT0 =  16'h69AA ;
    CCU2C addsub_6 (.A0(DataA[11]), .A1(DataA[12]), .B0(DataB[11]), .B1(DataB[12]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co5), 
        .S0(Result[11]), .S1(Result[12]), .COUT(co6));

    defparam addsub_7.INJECT1_1 = "NO" ;
    defparam addsub_7.INJECT1_0 = "NO" ;
    defparam addsub_7.INIT1 =  16'h69AA ;
    defparam addsub_7.INIT0 =  16'h69AA ;
    CCU2C addsub_7 (.A0(DataA[13]), .A1(DataA[14]), .B0(DataB[13]), .B1(DataB[14]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co6), 
        .S0(Result[13]), .S1(Result[14]), .COUT(co7));

    defparam addsub_8.INJECT1_1 = "NO" ;
    defparam addsub_8.INJECT1_0 = "NO" ;
    defparam addsub_8.INIT1 =  16'h69AA ;
    defparam addsub_8.INIT0 =  16'h69AA ;
    CCU2C addsub_8 (.A0(DataA[15]), .A1(DataA[16]), .B0(DataB[15]), .B1(DataB[16]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co7), 
        .S0(Result[15]), .S1(Result[16]), .COUT(co8));

    defparam addsub_9.INJECT1_1 = "NO" ;
    defparam addsub_9.INJECT1_0 = "NO" ;
    defparam addsub_9.INIT1 =  16'h69AA ;
    defparam addsub_9.INIT0 =  16'h69AA ;
    CCU2C addsub_9 (.A0(DataA[17]), .A1(DataA[18]), .B0(DataB[17]), .B1(DataB[18]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co8), 
        .S0(Result[17]), .S1(Result[18]), .COUT(co9));

    defparam addsub_10.INJECT1_1 = "NO" ;
    defparam addsub_10.INJECT1_0 = "NO" ;
    defparam addsub_10.INIT1 =  16'h69AA ;
    defparam addsub_10.INIT0 =  16'h69AA ;
    CCU2C addsub_10 (.A0(DataA[19]), .A1(DataA[20]), .B0(DataB[19]), .B1(DataB[20]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co9), 
        .S0(Result[19]), .S1(Result[20]), .COUT(co10));

    defparam addsub_11.INJECT1_1 = "NO" ;
    defparam addsub_11.INJECT1_0 = "NO" ;
    defparam addsub_11.INIT1 =  16'h69AA ;
    defparam addsub_11.INIT0 =  16'h69AA ;
    CCU2C addsub_11 (.A0(DataA[21]), .A1(DataA[22]), .B0(DataB[21]), .B1(DataB[22]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co10), 
        .S0(Result[21]), .S1(Result[22]), .COUT(co11));

    defparam addsub_12.INJECT1_1 = "NO" ;
    defparam addsub_12.INJECT1_0 = "NO" ;
    defparam addsub_12.INIT1 =  16'h69AA ;
    defparam addsub_12.INIT0 =  16'h69AA ;
    CCU2C addsub_12 (.A0(DataA[23]), .A1(DataA[24]), .B0(DataB[23]), .B1(DataB[24]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co11), 
        .S0(Result[23]), .S1(Result[24]), .COUT(co12));

    defparam addsub_13.INJECT1_1 = "NO" ;
    defparam addsub_13.INJECT1_0 = "NO" ;
    defparam addsub_13.INIT1 =  16'h69AA ;
    defparam addsub_13.INIT0 =  16'h69AA ;
    CCU2C addsub_13 (.A0(DataA[25]), .A1(DataA[26]), .B0(DataB[25]), .B1(DataB[26]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co12), 
        .S0(Result[25]), .S1(Result[26]), .COUT(co13));

    defparam addsub_14.INJECT1_1 = "NO" ;
    defparam addsub_14.INJECT1_0 = "NO" ;
    defparam addsub_14.INIT1 =  16'h69AA ;
    defparam addsub_14.INIT0 =  16'h69AA ;
    CCU2C addsub_14 (.A0(DataA[27]), .A1(DataA[28]), .B0(DataB[27]), .B1(DataB[28]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co13), 
        .S0(Result[27]), .S1(Result[28]), .COUT(co14));

    defparam addsub_15.INJECT1_1 = "NO" ;
    defparam addsub_15.INJECT1_0 = "NO" ;
    defparam addsub_15.INIT1 =  16'h69AA ;
    defparam addsub_15.INIT0 =  16'h69AA ;
    CCU2C addsub_15 (.A0(DataA[29]), .A1(DataA[30]), .B0(DataB[29]), .B1(DataB[30]), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co14), 
        .S0(Result[29]), .S1(Result[30]), .COUT(co15));

    defparam addsub_16.INJECT1_1 = "NO" ;
    defparam addsub_16.INJECT1_0 = "NO" ;
    defparam addsub_16.INIT1 =  16'h69AA ;
    defparam addsub_16.INIT0 =  16'h69AA ;
    CCU2C addsub_16 (.A0(DataA[31]), .A1(scuba_vlo), .B0(DataB[31]), .B1(add_sub_inv), 
        .C0(Add_Sub), .C1(Add_Sub), .D0(scuba_vhi), .D1(scuba_vhi), .CIN(co15), 
        .S0(Result[31]), .S1(Cout), .COUT(co16));

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam addsubd.INJECT1_1 = "NO" ;
    defparam addsubd.INJECT1_0 = "NO" ;
    defparam addsubd.INIT1 =  16'h66AA ;
    defparam addsubd.INIT0 =  16'h66AA ;
    CCU2C addsubd (.A0(scuba_vlo), .A1(scuba_vlo), .B0(scuba_vlo), .B1(scuba_vlo), 
        .C0(scuba_vhi), .C1(scuba_vhi), .D0(scuba_vhi), .D1(scuba_vhi), 
        .CIN(co16), .S0(co16d), .S1(), .COUT());



    // exemplar begin
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.12.1.454 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.12/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch sa5p00 -type bram -wp 10 -rp 0011 -data_width 1 -num_rows 32 -rdata_width 1 -read_reg1 outreg -gsr DISABLED -reset_rel async -memformat bin -cascade -1 -n pmi_ram_dpEbnonesadr153215321188cf97 -pmi -lang verilog  */
/* Sun Feb 06 15:10:23 2022 */


`timescale 1 ns / 1 ps
module pmi_ram_dpEbnonesadr153215321188cf97 (WrAddress, RdAddress, Data, 
    WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [4:0] WrAddress;
    input wire [4:0] RdAddress;
    input wire [0:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [0:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpEbnonesadr153215321188cf97_0_0_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr153215321188cf97_0_0_0.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr153215321188cf97_0_0_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr153215321188cf97_0_0_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr153215321188cf97_0_0_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr153215321188cf97_0_0_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr153215321188cf97_0_0_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr153215321188cf97_0_0_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr153215321188cf97_0_0_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr153215321188cf97_0_0_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr153215321188cf97_0_0_0.DATA_WIDTH_B = 1 ;
    defparam pmi_ram_dpEbnonesadr153215321188cf97_0_0_0.DATA_WIDTH_A = 1 ;
    DP16KD pmi_ram_dpEbnonesadr153215321188cf97_0_0_0 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), 
        .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), 
        .DIA0(Data[0]), .ADA13(scuba_vlo), .ADA12(scuba_vlo), .ADA11(scuba_vlo), 
        .ADA10(scuba_vlo), .ADA9(scuba_vlo), .ADA8(scuba_vlo), .ADA7(scuba_vlo), 
        .ADA6(scuba_vlo), .ADA5(scuba_vlo), .ADA4(WrAddress[4]), .ADA3(WrAddress[3]), 
        .ADA2(WrAddress[2]), .ADA1(WrAddress[1]), .ADA0(WrAddress[0]), .CEA(WrClockEn), 
        .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo), 
        .ADB13(scuba_vlo), .ADB12(scuba_vlo), .ADB11(scuba_vlo), .ADB10(scuba_vlo), 
        .ADB9(scuba_vlo), .ADB8(scuba_vlo), .ADB7(scuba_vlo), .ADB6(scuba_vlo), 
        .ADB5(scuba_vlo), .ADB4(RdAddress[4]), .ADB3(RdAddress[3]), .ADB2(RdAddress[2]), 
        .ADB1(RdAddress[1]), .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn), 
        .CLKB(RdClock), .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(Reset), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), 
        .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), 
        .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr153215321188cf97__PMIP__32__1__1B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpEbnonesadr153215321188cf97_0_0_0 MEM_LPC_FILE pmi_ram_dpEbnonesadr153215321188cf97__PMIP__32__1__1B
    // exemplar attribute pmi_ram_dpEbnonesadr153215321188cf97_0_0_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.12.1.454 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.12/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch sa5p00 -type bram -wp 10 -rp 0011 -data_width 150 -num_rows 2048 -rdata_width 150 -read_reg1 outreg -gsr DISABLED -reset_rel async -memformat bin -cascade -1 -n pmi_ram_dpEbnonesadr150112048150112048123cb5f0 -pmi -lang verilog  */
/* Sun Feb 06 15:10:23 2022 */


`timescale 1 ns / 1 ps
module pmi_ram_dpEbnonesadr150112048150112048123cb5f0 (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [10:0] WrAddress;
    input wire [10:0] RdAddress;
    input wire [149:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [149:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_0_16.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_0_16.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_0_16.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_0_16.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_0_16.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_0_16.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_0_16.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_0_16.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_0_16.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_0_16.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_0_16.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_0_16.DATA_WIDTH_A = 9 ;
    DP16KD pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_0_16 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(Data[8]), .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), 
        .DIA4(Data[4]), .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), 
        .DIA0(Data[0]), .ADA13(WrAddress[10]), .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), 
        .ADA10(WrAddress[7]), .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), 
        .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), 
        .ADA3(WrAddress[0]), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[10]), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), .DOA12(), .DOA11(), 
        .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), 
        .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), .DOB16(), .DOB15(), 
        .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(Q[8]), 
        .DOB7(Q[7]), .DOB6(Q[6]), .DOB5(Q[5]), .DOB4(Q[4]), .DOB3(Q[3]), 
        .DOB2(Q[2]), .DOB1(Q[1]), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_1_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_1_15.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_1_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_1_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_1_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_1_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_1_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_1_15.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_1_15.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_1_15.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_1_15.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_1_15.DATA_WIDTH_A = 9 ;
    DP16KD pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_1_15 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(Data[17]), .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), 
        .DIA4(Data[13]), .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), 
        .DIA0(Data[9]), .ADA13(WrAddress[10]), .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), 
        .ADA10(WrAddress[7]), .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), 
        .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), 
        .ADA3(WrAddress[0]), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[10]), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), .DOA12(), .DOA11(), 
        .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), 
        .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), .DOB16(), .DOB15(), 
        .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(Q[17]), 
        .DOB7(Q[16]), .DOB6(Q[15]), .DOB5(Q[14]), .DOB4(Q[13]), .DOB3(Q[12]), 
        .DOB2(Q[11]), .DOB1(Q[10]), .DOB0(Q[9]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_2_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_2_14.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_2_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_2_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_2_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_2_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_2_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_2_14.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_2_14.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_2_14.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_2_14.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_2_14.DATA_WIDTH_A = 9 ;
    DP16KD pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_2_14 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(Data[26]), .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), 
        .DIA4(Data[22]), .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), 
        .DIA0(Data[18]), .ADA13(WrAddress[10]), .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), 
        .ADA10(WrAddress[7]), .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), 
        .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), 
        .ADA3(WrAddress[0]), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[10]), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), .DOA12(), .DOA11(), 
        .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), 
        .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), .DOB16(), .DOB15(), 
        .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(Q[26]), 
        .DOB7(Q[25]), .DOB6(Q[24]), .DOB5(Q[23]), .DOB4(Q[22]), .DOB3(Q[21]), 
        .DOB2(Q[20]), .DOB1(Q[19]), .DOB0(Q[18]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_3_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_3_13.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_3_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_3_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_3_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_3_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_3_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_3_13.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_3_13.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_3_13.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_3_13.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_3_13.DATA_WIDTH_A = 9 ;
    DP16KD pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_3_13 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(Data[35]), .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), 
        .DIA4(Data[31]), .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), 
        .DIA0(Data[27]), .ADA13(WrAddress[10]), .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), 
        .ADA10(WrAddress[7]), .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), 
        .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), 
        .ADA3(WrAddress[0]), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[10]), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), .DOA12(), .DOA11(), 
        .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), 
        .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), .DOB16(), .DOB15(), 
        .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(Q[35]), 
        .DOB7(Q[34]), .DOB6(Q[33]), .DOB5(Q[32]), .DOB4(Q[31]), .DOB3(Q[30]), 
        .DOB2(Q[29]), .DOB1(Q[28]), .DOB0(Q[27]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_4_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_4_12.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_4_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_4_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_4_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_4_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_4_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_4_12.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_4_12.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_4_12.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_4_12.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_4_12.DATA_WIDTH_A = 9 ;
    DP16KD pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_4_12 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(Data[44]), .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), 
        .DIA4(Data[40]), .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), 
        .DIA0(Data[36]), .ADA13(WrAddress[10]), .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), 
        .ADA10(WrAddress[7]), .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), 
        .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), 
        .ADA3(WrAddress[0]), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[10]), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), .DOA12(), .DOA11(), 
        .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), 
        .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), .DOB16(), .DOB15(), 
        .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(Q[44]), 
        .DOB7(Q[43]), .DOB6(Q[42]), .DOB5(Q[41]), .DOB4(Q[40]), .DOB3(Q[39]), 
        .DOB2(Q[38]), .DOB1(Q[37]), .DOB0(Q[36]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_5_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_5_11.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_5_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_5_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_5_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_5_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_5_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_5_11.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_5_11.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_5_11.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_5_11.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_5_11.DATA_WIDTH_A = 9 ;
    DP16KD pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_5_11 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(Data[53]), .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), 
        .DIA4(Data[49]), .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), 
        .DIA0(Data[45]), .ADA13(WrAddress[10]), .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), 
        .ADA10(WrAddress[7]), .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), 
        .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), 
        .ADA3(WrAddress[0]), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[10]), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), .DOA12(), .DOA11(), 
        .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), 
        .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), .DOB16(), .DOB15(), 
        .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(Q[53]), 
        .DOB7(Q[52]), .DOB6(Q[51]), .DOB5(Q[50]), .DOB4(Q[49]), .DOB3(Q[48]), 
        .DOB2(Q[47]), .DOB1(Q[46]), .DOB0(Q[45]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_6_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_6_10.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_6_10.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_6_10.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_6_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_6_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_6_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_6_10.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_6_10.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_6_10.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_6_10.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_6_10.DATA_WIDTH_A = 9 ;
    DP16KD pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_6_10 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(Data[62]), .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), 
        .DIA4(Data[58]), .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), 
        .DIA0(Data[54]), .ADA13(WrAddress[10]), .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), 
        .ADA10(WrAddress[7]), .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), 
        .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), 
        .ADA3(WrAddress[0]), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[10]), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), .DOA12(), .DOA11(), 
        .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), 
        .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), .DOB16(), .DOB15(), 
        .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(Q[62]), 
        .DOB7(Q[61]), .DOB6(Q[60]), .DOB5(Q[59]), .DOB4(Q[58]), .DOB3(Q[57]), 
        .DOB2(Q[56]), .DOB1(Q[55]), .DOB0(Q[54]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_7_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_7_9.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_7_9.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_7_9.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_7_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_7_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_7_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_7_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_7_9.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_7_9.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_7_9.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_7_9.DATA_WIDTH_A = 9 ;
    DP16KD pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_7_9 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(Data[71]), .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), 
        .DIA4(Data[67]), .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), 
        .DIA0(Data[63]), .ADA13(WrAddress[10]), .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), 
        .ADA10(WrAddress[7]), .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), 
        .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), 
        .ADA3(WrAddress[0]), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[10]), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), .DOA12(), .DOA11(), 
        .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), 
        .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), .DOB16(), .DOB15(), 
        .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(Q[71]), 
        .DOB7(Q[70]), .DOB6(Q[69]), .DOB5(Q[68]), .DOB4(Q[67]), .DOB3(Q[66]), 
        .DOB2(Q[65]), .DOB1(Q[64]), .DOB0(Q[63]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_8_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_8_8.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_8_8.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_8_8.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_8_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_8_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_8_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_8_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_8_8.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_8_8.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_8_8.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_8_8.DATA_WIDTH_A = 9 ;
    DP16KD pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_8_8 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(Data[80]), .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), 
        .DIA4(Data[76]), .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), 
        .DIA0(Data[72]), .ADA13(WrAddress[10]), .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), 
        .ADA10(WrAddress[7]), .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), 
        .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), 
        .ADA3(WrAddress[0]), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[10]), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), .DOA12(), .DOA11(), 
        .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), 
        .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), .DOB16(), .DOB15(), 
        .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(Q[80]), 
        .DOB7(Q[79]), .DOB6(Q[78]), .DOB5(Q[77]), .DOB4(Q[76]), .DOB3(Q[75]), 
        .DOB2(Q[74]), .DOB1(Q[73]), .DOB0(Q[72]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_9_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_9_7.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_9_7.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_9_7.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_9_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_9_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_9_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_9_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_9_7.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_9_7.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_9_7.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_9_7.DATA_WIDTH_A = 9 ;
    DP16KD pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_9_7 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(Data[89]), .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), 
        .DIA4(Data[85]), .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), 
        .DIA0(Data[81]), .ADA13(WrAddress[10]), .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), 
        .ADA10(WrAddress[7]), .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), 
        .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), 
        .ADA3(WrAddress[0]), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[10]), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), .DOA12(), .DOA11(), 
        .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), 
        .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), .DOB16(), .DOB15(), 
        .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(Q[89]), 
        .DOB7(Q[88]), .DOB6(Q[87]), .DOB5(Q[86]), .DOB4(Q[85]), .DOB3(Q[84]), 
        .DOB2(Q[83]), .DOB1(Q[82]), .DOB0(Q[81]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_10_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_10_6.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_10_6.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_10_6.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_10_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_10_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_10_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_10_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_10_6.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_10_6.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_10_6.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_10_6.DATA_WIDTH_A = 9 ;
    DP16KD pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_10_6 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(Data[98]), .DIA7(Data[97]), .DIA6(Data[96]), .DIA5(Data[95]), 
        .DIA4(Data[94]), .DIA3(Data[93]), .DIA2(Data[92]), .DIA1(Data[91]), 
        .DIA0(Data[90]), .ADA13(WrAddress[10]), .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), 
        .ADA10(WrAddress[7]), .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), 
        .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), 
        .ADA3(WrAddress[0]), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[10]), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), .DOA12(), .DOA11(), 
        .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), 
        .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), .DOB16(), .DOB15(), 
        .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(Q[98]), 
        .DOB7(Q[97]), .DOB6(Q[96]), .DOB5(Q[95]), .DOB4(Q[94]), .DOB3(Q[93]), 
        .DOB2(Q[92]), .DOB1(Q[91]), .DOB0(Q[90]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_11_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_11_5.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_11_5.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_11_5.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_11_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_11_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_11_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_11_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_11_5.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_11_5.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_11_5.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_11_5.DATA_WIDTH_A = 9 ;
    DP16KD pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_11_5 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(Data[107]), .DIA7(Data[106]), .DIA6(Data[105]), .DIA5(Data[104]), 
        .DIA4(Data[103]), .DIA3(Data[102]), .DIA2(Data[101]), .DIA1(Data[100]), 
        .DIA0(Data[99]), .ADA13(WrAddress[10]), .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), 
        .ADA10(WrAddress[7]), .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), 
        .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), 
        .ADA3(WrAddress[0]), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[10]), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), .DOA12(), .DOA11(), 
        .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), 
        .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), .DOB16(), .DOB15(), 
        .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(Q[107]), 
        .DOB7(Q[106]), .DOB6(Q[105]), .DOB5(Q[104]), .DOB4(Q[103]), .DOB3(Q[102]), 
        .DOB2(Q[101]), .DOB1(Q[100]), .DOB0(Q[99]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_12_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_12_4.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_12_4.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_12_4.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_12_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_12_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_12_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_12_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_12_4.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_12_4.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_12_4.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_12_4.DATA_WIDTH_A = 9 ;
    DP16KD pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_12_4 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(Data[116]), .DIA7(Data[115]), .DIA6(Data[114]), .DIA5(Data[113]), 
        .DIA4(Data[112]), .DIA3(Data[111]), .DIA2(Data[110]), .DIA1(Data[109]), 
        .DIA0(Data[108]), .ADA13(WrAddress[10]), .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), 
        .ADA10(WrAddress[7]), .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), 
        .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), 
        .ADA3(WrAddress[0]), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[10]), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), .DOA12(), .DOA11(), 
        .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), 
        .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), .DOB16(), .DOB15(), 
        .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(Q[116]), 
        .DOB7(Q[115]), .DOB6(Q[114]), .DOB5(Q[113]), .DOB4(Q[112]), .DOB3(Q[111]), 
        .DOB2(Q[110]), .DOB1(Q[109]), .DOB0(Q[108]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_13_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_13_3.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_13_3.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_13_3.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_13_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_13_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_13_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_13_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_13_3.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_13_3.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_13_3.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_13_3.DATA_WIDTH_A = 9 ;
    DP16KD pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_13_3 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(Data[125]), .DIA7(Data[124]), .DIA6(Data[123]), .DIA5(Data[122]), 
        .DIA4(Data[121]), .DIA3(Data[120]), .DIA2(Data[119]), .DIA1(Data[118]), 
        .DIA0(Data[117]), .ADA13(WrAddress[10]), .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), 
        .ADA10(WrAddress[7]), .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), 
        .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), 
        .ADA3(WrAddress[0]), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[10]), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), .DOA12(), .DOA11(), 
        .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), 
        .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), .DOB16(), .DOB15(), 
        .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(Q[125]), 
        .DOB7(Q[124]), .DOB6(Q[123]), .DOB5(Q[122]), .DOB4(Q[121]), .DOB3(Q[120]), 
        .DOB2(Q[119]), .DOB1(Q[118]), .DOB0(Q[117]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_14_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_14_2.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_14_2.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_14_2.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_14_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_14_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_14_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_14_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_14_2.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_14_2.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_14_2.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_14_2.DATA_WIDTH_A = 9 ;
    DP16KD pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_14_2 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(Data[134]), .DIA7(Data[133]), .DIA6(Data[132]), .DIA5(Data[131]), 
        .DIA4(Data[130]), .DIA3(Data[129]), .DIA2(Data[128]), .DIA1(Data[127]), 
        .DIA0(Data[126]), .ADA13(WrAddress[10]), .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), 
        .ADA10(WrAddress[7]), .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), 
        .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), 
        .ADA3(WrAddress[0]), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[10]), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), .DOA12(), .DOA11(), 
        .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), 
        .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), .DOB16(), .DOB15(), 
        .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(Q[134]), 
        .DOB7(Q[133]), .DOB6(Q[132]), .DOB5(Q[131]), .DOB4(Q[130]), .DOB3(Q[129]), 
        .DOB2(Q[128]), .DOB1(Q[127]), .DOB0(Q[126]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_15_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_15_1.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_15_1.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_15_1.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_15_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_15_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_15_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_15_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_15_1.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_15_1.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_15_1.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_15_1.DATA_WIDTH_A = 9 ;
    DP16KD pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_15_1 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(Data[143]), .DIA7(Data[142]), .DIA6(Data[141]), .DIA5(Data[140]), 
        .DIA4(Data[139]), .DIA3(Data[138]), .DIA2(Data[137]), .DIA1(Data[136]), 
        .DIA0(Data[135]), .ADA13(WrAddress[10]), .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), 
        .ADA10(WrAddress[7]), .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), 
        .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), 
        .ADA3(WrAddress[0]), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[10]), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), .DOA12(), .DOA11(), 
        .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), 
        .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), .DOB16(), .DOB15(), 
        .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(Q[143]), 
        .DOB7(Q[142]), .DOB6(Q[141]), .DOB5(Q[140]), .DOB4(Q[139]), .DOB3(Q[138]), 
        .DOB2(Q[137]), .DOB1(Q[136]), .DOB0(Q[135]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B" */
             /* synthesis MEM_INIT_FILE="" */;

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_16_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_16_0.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_16_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_16_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_16_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_16_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_16_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_16_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_16_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_16_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_16_0.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_16_0.DATA_WIDTH_A = 9 ;
    DP16KD pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_16_0 (.DIA17(scuba_vlo), 
        .DIA16(scuba_vlo), .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), 
        .DIA12(scuba_vlo), .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), 
        .DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(Data[149]), 
        .DIA4(Data[148]), .DIA3(Data[147]), .DIA2(Data[146]), .DIA1(Data[145]), 
        .DIA0(Data[144]), .ADA13(WrAddress[10]), .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), 
        .ADA10(WrAddress[7]), .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), 
        .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), 
        .ADA3(WrAddress[0]), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB17(scuba_vlo), 
        .DIB16(scuba_vlo), .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), 
        .DIB12(scuba_vlo), .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), 
        .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), 
        .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), 
        .DIB0(scuba_vlo), .ADB13(RdAddress[10]), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(Reset), 
        .DOA17(), .DOA16(), .DOA15(), .DOA14(), .DOA13(), .DOA12(), .DOA11(), 
        .DOA10(), .DOA9(), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), 
        .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB17(), .DOB16(), .DOB15(), 
        .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(), 
        .DOB7(), .DOB6(), .DOB5(Q[149]), .DOB4(Q[148]), .DOB3(Q[147]), .DOB2(Q[146]), 
        .DOB1(Q[145]), .DOB0(Q[144]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_0_16 MEM_LPC_FILE pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_0_16 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_1_15 MEM_LPC_FILE pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_1_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_2_14 MEM_LPC_FILE pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_2_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_3_13 MEM_LPC_FILE pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_3_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_4_12 MEM_LPC_FILE pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_4_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_5_11 MEM_LPC_FILE pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_5_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_6_10 MEM_LPC_FILE pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_6_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_7_9 MEM_LPC_FILE pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_7_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_8_8 MEM_LPC_FILE pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_8_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_9_7 MEM_LPC_FILE pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_9_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_10_6 MEM_LPC_FILE pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_10_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_11_5 MEM_LPC_FILE pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_11_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_12_4 MEM_LPC_FILE pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_12_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_13_3 MEM_LPC_FILE pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_13_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_14_2 MEM_LPC_FILE pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_14_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_15_1 MEM_LPC_FILE pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_15_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_16_0 MEM_LPC_FILE pmi_ram_dpEbnonesadr150112048150112048123cb5f0__PMIP__2048__150__150B
    // exemplar attribute pmi_ram_dpEbnonesadr150112048150112048123cb5f0_0_16_0 MEM_INIT_FILE 
    // exemplar end

endmodule
